// *************************************************************
// Created by David J. Marion aka FPGA Dude
// A ROM containing patterns for ASCII values.
//
// Non-printable characters 00 - 1f, and 7f
// Printable characters 20 - 7e
//
// Not all character ROMs have been patterned.
// Only numbers, capital letters, some spec chars. 
//		Numbers       30 - 39
//   	Letters       41 - 5a 
//      (smiley face)   01
//		(space)         20
//		   .            2e
// 		   :            3a
//		   |	        7c	
//
// The 7-bit ASCII code for each character is used as
// the MSB of the address. The 4-bit LSB is the row value.
// *************************************************************

module ascii_rom(
	input clk, 
	input wire [15:0] addr,
	output reg [7:0] data
	);

	(* rom_style = "block" *)	// Infer BRAM

	reg [15:0] addr_reg;
	
	always @(posedge clk)
		addr_reg <= addr;
		
	always @*
		case(addr_reg)
			// Begin non-printable ASCII characters (00 - 1f)
			// code x0000 (nul) null byte, which is the all-zero pattern
			16'h0000: data = 8'b00000000;	//
			16'h0001: data = 8'b00000000;	//
			16'h0002: data = 8'b00000000;	//
			16'h0003: data = 8'b00000000;	//
			16'h0004: data = 8'b00000000;	//
			16'h0005: data = 8'b00000000;	//
			16'h0006: data = 8'b00000000;	//
			16'h0007: data = 8'b00000000;	//
			16'h0008: data = 8'b00000000;	//
			16'h0009: data = 8'b00000000;	//
			16'h000a: data = 8'b00000000;	//
			16'h000b: data = 8'b00000000;	//
			16'h000c: data = 8'b00000000;	//
			16'h000d: data = 8'b00000000;	//
			16'h000e: data = 8'b00000000;	//
			16'h000f: data = 8'b00000000;	//
			// code x0001 (soh) start of heading
			16'h0010: data = 8'b00000000;	//
			16'h0011: data = 8'b00000000;	//
			16'h0012: data = 8'b01111110;	// ******			
			16'h0013: data = 8'b10000001;	//*      *
			16'h0014: data = 8'b10100101;	//* *  * *
			16'h0015: data = 8'b10000001;	//*      *
			16'h0016: data = 8'b10000001;	//*      *
			16'h0017: data = 8'b10111101;	//* **** *
			16'h0018: data = 8'b10011001;	//*  **  *
			16'h0019: data = 8'b10000001;	//*      *
			16'h001a: data = 8'b10000001;	//*      *
			16'h001b: data = 8'b01111110;	// ******
			16'h001c: data = 8'b00000000;	//
			16'h001d: data = 8'b00000000;	//
			16'h001e: data = 8'b00000000;	//
			16'h001f: data = 8'b00000000;	//
			// code x0002 (stx) start of text
			16'h0020: data = 8'b00000000;	//
			16'h0021: data = 8'b00000000;	//
			16'h0022: data = 8'b00000000;	//
			16'h0023: data = 8'b00000000;	//
			16'h0024: data = 8'b00000000;	//
			16'h0025: data = 8'b00000000;	//
			16'h0026: data = 8'b00000000;	//
			16'h0027: data = 8'b00000000;	//
			16'h0028: data = 8'b00000000;	//
			16'h0029: data = 8'b00000000;	//
			16'h002a: data = 8'b00000000;	//
			16'h002b: data = 8'b00000000;	//
			16'h002c: data = 8'b00000000;	//
			16'h002d: data = 8'b00000000;	//
			16'h002e: data = 8'b00000000;	//
			16'h002f: data = 8'b00000000;	//
			// code x0003 (etx) end of text
			16'h0030: data = 8'b00000000;	//
			16'h0031: data = 8'b00000000;	//
			16'h0032: data = 8'b00000000;	//
			16'h0033: data = 8'b00000000;	//
			16'h0034: data = 8'b00000000;	//
			16'h0035: data = 8'b00000000;	//
			16'h0036: data = 8'b00000000;	//
			16'h0037: data = 8'b00000000;	//
			16'h0038: data = 8'b00000000;	//
			16'h0039: data = 8'b00000000;	//
			16'h003a: data = 8'b00000000;	//
			16'h003b: data = 8'b00000000;	//
			16'h003c: data = 8'b00000000;	//
			16'h003d: data = 8'b00000000;	//
			16'h003e: data = 8'b00000000;	//
			16'h003f: data = 8'b00000000;	//
			// code x0004 (eot) end of transmission
			16'h0040: data = 8'b00000000;	//
			16'h0041: data = 8'b00000000;	//
			16'h0042: data = 8'b00000000;	//
			16'h0043: data = 8'b00000000;	//
			16'h0044: data = 8'b00000000;	//
			16'h0045: data = 8'b00000000;	//
			16'h0046: data = 8'b00000000;	//
			16'h0047: data = 8'b00000000;	//
			16'h0048: data = 8'b00000000;	//
			16'h0049: data = 8'b00000000;	//
			16'h004a: data = 8'b00000000;	//
			16'h004b: data = 8'b00000000;	//
			16'h004c: data = 8'b00000000;	//
			16'h004d: data = 8'b00000000;	//
			16'h004e: data = 8'b00000000;	//
			16'h004f: data = 8'b00000000;	//
			// code x0005 (enq) end of query
			16'h0050: data = 8'b00000000;	//
			16'h0051: data = 8'b00000000;	//
			16'h0052: data = 8'b00000000;	//
			16'h0053: data = 8'b00000000;	//
			16'h0054: data = 8'b00000000;	//
			16'h0055: data = 8'b00000000;	//
			16'h0056: data = 8'b00000000;	//
			16'h0057: data = 8'b00000000;	//
			16'h0058: data = 8'b00000000;	//
			16'h0059: data = 8'b00000000;	//
			16'h005a: data = 8'b00000000;	//
			16'h005b: data = 8'b00000000;	//
			16'h005c: data = 8'b00000000;	//
			16'h005d: data = 8'b00000000;	//
			16'h005e: data = 8'b00000000;	//
			16'h005f: data = 8'b00000000;	//
			// code x0006 (ack) acknowledge
			16'h0060: data = 8'b00000000;	//
			16'h0061: data = 8'b00000000;	//
			16'h0062: data = 8'b00000000;	//
			16'h0063: data = 8'b00000000;	//
			16'h0064: data = 8'b00000000;	//
			16'h0065: data = 8'b00000000;	//
			16'h0066: data = 8'b00000000;	//
			16'h0067: data = 8'b00000000;	//
			16'h0068: data = 8'b00000000;	//
			16'h0069: data = 8'b00000000;	//
			16'h006a: data = 8'b00000000;	//
			16'h006b: data = 8'b00000000;	//
			16'h006c: data = 8'b00000000;	//
			16'h006d: data = 8'b00000000;	//
			16'h006e: data = 8'b00000000;	//
			16'h006f: data = 8'b00000000;	//
			// code x0007 (bel) generate a bell sound, if supported
			16'h0070: data = 8'b00000000;	//
			16'h0071: data = 8'b00000000;	//
			16'h0072: data = 8'b00000000;	//
			16'h0073: data = 8'b00000000;	//
			16'h0074: data = 8'b00000000;	//
			16'h0075: data = 8'b00000000;	//
			16'h0076: data = 8'b00000000;	//
			16'h0077: data = 8'b00000000;	//
			16'h0078: data = 8'b00000000;	//
			16'h0079: data = 8'b00000000;	//
			16'h007a: data = 8'b00000000;	//
			16'h007b: data = 8'b00000000;	//
			16'h007c: data = 8'b00000000;	//
			16'h007d: data = 8'b00000000;	//
			16'h007e: data = 8'b00000000;	//
			16'h007f: data = 8'b00000000;	//
			// code x0008 (bs) backspace
			16'h0080: data = 8'b00000000;	//
			16'h0081: data = 8'b00000000;	//
			16'h0082: data = 8'b00000000;	//
			16'h0083: data = 8'b00000000;	//
			16'h0084: data = 8'b00000000;	//
			16'h0085: data = 8'b00000000;	//
			16'h0086: data = 8'b00000000;	//
			16'h0087: data = 8'b00000000;	//
			16'h0088: data = 8'b00000000;	//
			16'h0089: data = 8'b00000000;	//
			16'h008a: data = 8'b00000000;	//
			16'h008b: data = 8'b00000000;	//
			16'h008c: data = 8'b00000000;	//
			16'h008d: data = 8'b00000000;	//
			16'h008e: data = 8'b00000000;	//
			16'h008f: data = 8'b00000000;	//
			// code x0009 (ht) horizontal tab
			16'h0090: data = 8'b00000000;	//
			16'h0091: data = 8'b00000000;	//
			16'h0092: data = 8'b00000000;	//
			16'h0093: data = 8'b00000000;	//
			16'h0094: data = 8'b00000000;	//
			16'h0095: data = 8'b00000000;	//
			16'h0096: data = 8'b00000000;	//
			16'h0097: data = 8'b00000000;	//
			16'h0098: data = 8'b00000000;	//
			16'h0099: data = 8'b00000000;	//
			16'h009a: data = 8'b00000000;	//
			16'h009b: data = 8'b00000000;	//
			16'h009c: data = 8'b00000000;	//
			16'h009d: data = 8'b00000000;	//
			16'h009e: data = 8'b00000000;	//
			16'h009f: data = 8'b00000000;	//
			// code x000a (nl) new line
			16'h00a0: data = 8'b00000000;	//
			16'h00a1: data = 8'b00000000;	//
			16'h00a2: data = 8'b00000000;	//
			16'h00a3: data = 8'b00000000;	//
			16'h00a4: data = 8'b00000000;	//
			16'h00a5: data = 8'b00000000;	//
			16'h00a6: data = 8'b00000000;	//
			16'h00a7: data = 8'b00000000;	//
			16'h00a8: data = 8'b00000000;	//
			16'h00a9: data = 8'b00000000;	//
			16'h00aa: data = 8'b00000000;	//
			16'h00ab: data = 8'b00000000;	//
			16'h00ac: data = 8'b00000000;	//
			16'h00ad: data = 8'b00000000;	//
			16'h00ae: data = 8'b00000000;	//
			16'h00af: data = 8'b00000000;	//
			// code x000b (vt) vertical tab
			16'h00b0: data = 8'b00000000;	//
			16'h00b1: data = 8'b00000000;	//
			16'h00b2: data = 8'b00000000;	//
			16'h00b3: data = 8'b00000000;	//
			16'h00b4: data = 8'b00000000;	//
			16'h00b5: data = 8'b00000000;	//
			16'h00b6: data = 8'b00000000;	//
			16'h00b7: data = 8'b00000000;	//
			16'h00b8: data = 8'b00000000;	//
			16'h00b9: data = 8'b00000000;	//
			16'h00ba: data = 8'b00000000;	//
			16'h00bb: data = 8'b00000000;	//
			16'h00bc: data = 8'b00000000;	//
			16'h00bd: data = 8'b00000000;	//
			16'h00be: data = 8'b00000000;	//
			16'h00bf: data = 8'b00000000;	//
			// code x000c (np) new page
			16'h00c0: data = 8'b00000000;	//
			16'h00c1: data = 8'b00000000;	//
			16'h00c2: data = 8'b00000000;	//
			16'h00c3: data = 8'b00000000;	//
			16'h00c4: data = 8'b00000000;	//
			16'h00c5: data = 8'b00000000;	//
			16'h00c6: data = 8'b00000000;	//
			16'h00c7: data = 8'b00000000;	//
			16'h00c8: data = 8'b00000000;	//
			16'h00c9: data = 8'b00000000;	//
			16'h00ca: data = 8'b00000000;	//
			16'h00cb: data = 8'b00000000;	//
			16'h00cc: data = 8'b00000000;	//
			16'h00cd: data = 8'b00000000;	//
			16'h00ce: data = 8'b00000000;	//
			16'h00cf: data = 8'b00000000;	//
			// code x000d (cr) carriage return
			16'h00d0: data = 8'b00000000;	//
			16'h00d1: data = 8'b00000000;	//
			16'h00d2: data = 8'b00000000;	//
			16'h00d3: data = 8'b00000000;	//
			16'h00d4: data = 8'b00000000;	//
			16'h00d5: data = 8'b00000000;	//
			16'h00d6: data = 8'b00000000;	//
			16'h00d7: data = 8'b00000000;	//
			16'h00d8: data = 8'b00000000;	//
			16'h00d9: data = 8'b00000000;	//
			16'h00da: data = 8'b00000000;	//
			16'h00db: data = 8'b00000000;	//
			16'h00dc: data = 8'b00000000;	//
			16'h00dd: data = 8'b00000000;	//
			16'h00de: data = 8'b00000000;	//
			16'h00df: data = 8'b00000000;	//
			// code x000e (so) shift out
			16'h00e0: data = 8'b00000000;	//
			16'h00e1: data = 8'b00000000;	//
			16'h00e2: data = 8'b00000000;	//
			16'h00e3: data = 8'b00000000;	//
			16'h00e4: data = 8'b00000000;	//
			16'h00e5: data = 8'b00000000;	//
			16'h00e6: data = 8'b00000000;	//
			16'h00e7: data = 8'b00000000;	//
			16'h00e8: data = 8'b00000000;	//
			16'h00e9: data = 8'b00000000;	//
			16'h00ea: data = 8'b00000000;	//
			16'h00eb: data = 8'b00000000;	//
			16'h00ec: data = 8'b00000000;	//
			16'h00ed: data = 8'b00000000;	//
			16'h00ee: data = 8'b00000000;	//
			16'h00ef: data = 8'b00000000;	//
			// code x000f (si) shift in
			16'h00f0: data = 8'b00000000;	//
			16'h00f1: data = 8'b00000000;	//
			16'h00f2: data = 8'b00000000;	//
			16'h00f3: data = 8'b00000000;	//
			16'h00f4: data = 8'b00000000;	//
			16'h00f5: data = 8'b00000000;	//
			16'h00f6: data = 8'b00000000;	//
			16'h00f7: data = 8'b00000000;	//
			16'h00f8: data = 8'b00000000;	//
			16'h00f9: data = 8'b00000000;	//
			16'h00fa: data = 8'b00000000;	//
			16'h00fb: data = 8'b00000000;	//
			16'h00fc: data = 8'b00000000;	//
			16'h00fd: data = 8'b00000000;	//
			16'h00fe: data = 8'b00000000;	//
			16'h00ff: data = 8'b00000000;	//
			// code x0010 (dle) data link escape
			16'h0100: data = 8'b00000000;	//
			16'h0101: data = 8'b00000000;	//
			16'h0102: data = 8'b00000000;	//
			16'h0103: data = 8'b00000000;	//
			16'h0104: data = 8'b00000000;	//
			16'h0105: data = 8'b00000000;	//
			16'h0106: data = 8'b00000000;	//
			16'h0107: data = 8'b00000000;	//
			16'h0108: data = 8'b00000000;	//
			16'h0109: data = 8'b00000000;	//
			16'h010a: data = 8'b00000000;	//
			16'h010b: data = 8'b00000000;	//
			16'h010c: data = 8'b00000000;	//
			16'h010d: data = 8'b00000000;	//
			16'h010e: data = 8'b00000000;	//
			16'h010f: data = 8'b00000000;	//
			// code x0011 (dc1) device control 1
			16'h0110: data = 8'b00000000;	//
			16'h0111: data = 8'b00000000;	//
			16'h0112: data = 8'b00000000;	//
			16'h0113: data = 8'b00000000;	//
			16'h0114: data = 8'b00000000;	//
			16'h0115: data = 8'b00000000;	//
			16'h0116: data = 8'b00000000;	//
			16'h0117: data = 8'b00000000;	//
			16'h0118: data = 8'b00000000;	//
			16'h0119: data = 8'b00000000;	//
			16'h011a: data = 8'b00000000;	//
			16'h011b: data = 8'b00000000;	//
			16'h011c: data = 8'b00000000;	//
			16'h011d: data = 8'b00000000;	//
			16'h011e: data = 8'b00000000;	//
			16'h011f: data = 8'b00000000;	//
			// code x0012 (dc2) device control 2
			16'h0120: data = 8'b00000000;	//
			16'h0121: data = 8'b00000000;	//
			16'h0122: data = 8'b00000000;	//
			16'h0123: data = 8'b00000000;	//
			16'h0124: data = 8'b00000000;	//
			16'h0125: data = 8'b00000000;	//
			16'h0126: data = 8'b00000000;	//
			16'h0127: data = 8'b00000000;	//
			16'h0128: data = 8'b00000000;	//
			16'h0129: data = 8'b00000000;	//
			16'h012a: data = 8'b00000000;	//
			16'h012b: data = 8'b00000000;	//
			16'h012c: data = 8'b00000000;	//
			16'h012d: data = 8'b00000000;	//
			16'h012e: data = 8'b00000000;	//
			16'h012f: data = 8'b00000000;	//
			// code x0013 (dc3) device control 3
			16'h0130: data = 8'b00000000;	//
			16'h0131: data = 8'b00000000;	//
			16'h0132: data = 8'b00000000;	//
			16'h0133: data = 8'b00000000;	//
			16'h0134: data = 8'b00000000;	//
			16'h0135: data = 8'b00000000;	//
			16'h0136: data = 8'b00000000;	//
			16'h0137: data = 8'b00000000;	//
			16'h0138: data = 8'b00000000;	//
			16'h0139: data = 8'b00000000;	//
			16'h013a: data = 8'b00000000;	//
			16'h013b: data = 8'b00000000;	//
			16'h013c: data = 8'b00000000;	//
			16'h013d: data = 8'b00000000;	//
			16'h013e: data = 8'b00000000;	//
			16'h013f: data = 8'b00000000;	//
			// code x0014 (dc4) device control 4
			16'h0140: data = 8'b00000000;	//
			16'h0141: data = 8'b00000000;	//
			16'h0142: data = 8'b00000000;	//
			16'h0143: data = 8'b00000000;	//
			16'h0144: data = 8'b00000000;	//
			16'h0145: data = 8'b00000000;	//
			16'h0146: data = 8'b00000000;	//
			16'h0147: data = 8'b00000000;	//
			16'h0148: data = 8'b00000000;	//
			16'h0149: data = 8'b00000000;	//
			16'h014a: data = 8'b00000000;	//
			16'h014b: data = 8'b00000000;	//
			16'h014c: data = 8'b00000000;	//
			16'h014d: data = 8'b00000000;	//
			16'h014e: data = 8'b00000000;	//
			16'h014f: data = 8'b00000000;	//
			// code x0015 (nak) negative acknowledgement
			16'h0150: data = 8'b00000000;	//
			16'h0151: data = 8'b00000000;	//
			16'h0152: data = 8'b00000000;	//
			16'h0153: data = 8'b00000000;	//
			16'h0154: data = 8'b00000000;	//
			16'h0155: data = 8'b00000000;	//
			16'h0156: data = 8'b00000000;	//
			16'h0157: data = 8'b00000000;	//
			16'h0158: data = 8'b00000000;	//
			16'h0159: data = 8'b00000000;	//
			16'h015a: data = 8'b00000000;	//
			16'h015b: data = 8'b00000000;	//
			16'h015c: data = 8'b00000000;	//
			16'h015d: data = 8'b00000000;	//
			16'h015e: data = 8'b00000000;	//
			16'h015f: data = 8'b00000000;	//
			// code x0016 (syn) synchronize
			16'h0160: data = 8'b00000000;	//
			16'h0161: data = 8'b00000000;	//
			16'h0162: data = 8'b00000000;	//
			16'h0163: data = 8'b00000000;	//
			16'h0164: data = 8'b00000000;	//
			16'h0165: data = 8'b00000000;	//
			16'h0166: data = 8'b00000000;	//
			16'h0167: data = 8'b00000000;	//
			16'h0168: data = 8'b00000000;	//
			16'h0169: data = 8'b00000000;	//
			16'h016a: data = 8'b00000000;	//
			16'h016b: data = 8'b00000000;	//
			16'h016c: data = 8'b00000000;	//
			16'h016d: data = 8'b00000000;	//
			16'h016e: data = 8'b00000000;	//
			16'h016f: data = 8'b00000000;	//
			// code x0017 (etb) end of transmission block
			16'h0170: data = 8'b00000000;	//
			16'h0171: data = 8'b00000000;	//
			16'h0172: data = 8'b00000000;	//
			16'h0173: data = 8'b00000000;	//
			16'h0174: data = 8'b00000000;	//
			16'h0175: data = 8'b00000000;	//
			16'h0176: data = 8'b00000000;	//
			16'h0177: data = 8'b00000000;	//
			16'h0178: data = 8'b00000000;	//
			16'h0179: data = 8'b00000000;	//
			16'h017a: data = 8'b00000000;	//
			16'h017b: data = 8'b00000000;	//
			16'h017c: data = 8'b00000000;	//
			16'h017d: data = 8'b00000000;	//
			16'h017e: data = 8'b00000000;	//
			16'h017f: data = 8'b00000000;	//
			// code x0018 (can) cancel
			16'h0180: data = 8'b00000000;	//
			16'h0181: data = 8'b00000000;	//
			16'h0182: data = 8'b00000000;	//
			16'h0183: data = 8'b00000000;	//
			16'h0184: data = 8'b00000000;	//
			16'h0185: data = 8'b00000000;	//
			16'h0186: data = 8'b00000000;	//
			16'h0187: data = 8'b00000000;	//
			16'h0188: data = 8'b00000000;	//
			16'h0189: data = 8'b00000000;	//
			16'h018a: data = 8'b00000000;	//
			16'h018b: data = 8'b00000000;	//
			16'h018c: data = 8'b00000000;	//
			16'h018d: data = 8'b00000000;	//
			16'h018e: data = 8'b00000000;	//
			16'h018f: data = 8'b00000000;	//
			// code x0019 (em) end of medium
			16'h0190: data = 8'b00000000;	//
			16'h0191: data = 8'b00000000;	//
			16'h0192: data = 8'b00000000;	//
			16'h0193: data = 8'b00000000;	//
			16'h0194: data = 8'b00000000;	//
			16'h0195: data = 8'b00000000;	//
			16'h0196: data = 8'b00000000;	//
			16'h0197: data = 8'b00000000;	//
			16'h0198: data = 8'b00000000;	//
			16'h0199: data = 8'b00000000;	//
			16'h019a: data = 8'b00000000;	//
			16'h019b: data = 8'b00000000;	//
			16'h019c: data = 8'b00000000;	//
			16'h019d: data = 8'b00000000;	//
			16'h019e: data = 8'b00000000;	//
			16'h019f: data = 8'b00000000;	//
			// code x001a (sub) substitute
			16'h01a0: data = 8'b00000000;	//
			16'h01a1: data = 8'b00000000;	//
			16'h01a2: data = 8'b00000000;	//
			16'h01a3: data = 8'b00000000;	//
			16'h01a4: data = 8'b00000000;	//
			16'h01a5: data = 8'b00000000;	//
			16'h01a6: data = 8'b00000000;	//
			16'h01a7: data = 8'b00000000;	//
			16'h01a8: data = 8'b00000000;	//
			16'h01a9: data = 8'b00000000;	//
			16'h01aa: data = 8'b00000000;	//
			16'h01ab: data = 8'b00000000;	//
			16'h01ac: data = 8'b00000000;	//
			16'h01ad: data = 8'b00000000;	//
			16'h01ae: data = 8'b00000000;	//
			16'h01af: data = 8'b00000000;	//
			// code x001b (esc) escape
			16'h01b0: data = 8'b00000000;	//
			16'h01b1: data = 8'b00000000;	//
			16'h01b2: data = 8'b00000000;	//
			16'h01b3: data = 8'b00000000;	//
			16'h01b4: data = 8'b00000000;	//
			16'h01b5: data = 8'b00000000;	//
			16'h01b6: data = 8'b00000000;	//
			16'h01b7: data = 8'b00000000;	//
			16'h01b8: data = 8'b00000000;	//
			16'h01b9: data = 8'b00000000;	//
			16'h01ba: data = 8'b00000000;	//
			16'h01bb: data = 8'b00000000;	//
			16'h01bc: data = 8'b00000000;	//
			16'h01bd: data = 8'b00000000;	//
			16'h01be: data = 8'b00000000;	//
			16'h01bf: data = 8'b00000000;	//
			// code x001c (fs) file separator
			16'h01c0: data = 8'b00000000;	//
			16'h01c1: data = 8'b00000000;	//
			16'h01c2: data = 8'b00000000;	//
			16'h01c3: data = 8'b00000000;	//
			16'h01c4: data = 8'b00000000;	//
			16'h01c5: data = 8'b00000000;	//
			16'h01c6: data = 8'b00000000;	//
			16'h01c7: data = 8'b00000000;	//
			16'h01c8: data = 8'b00000000;	//
			16'h01c9: data = 8'b00000000;	//
			16'h01ca: data = 8'b00000000;	//
			16'h01cb: data = 8'b00000000;	//
			16'h01cc: data = 8'b00000000;	//
			16'h01cd: data = 8'b00000000;	//
			16'h01ce: data = 8'b00000000;	//
			16'h01cf: data = 8'b00000000;	//
			// code x001d (gs) group separator
			16'h01d0: data = 8'b00000000;	//
			16'h01d1: data = 8'b00000000;	//
			16'h01d2: data = 8'b00000000;	//
			16'h01d3: data = 8'b00000000;	//
			16'h01d4: data = 8'b00000000;	//
			16'h01d5: data = 8'b00000000;	//
			16'h01d6: data = 8'b00000000;	//
			16'h01d7: data = 8'b00000000;	//
			16'h01d8: data = 8'b00000000;	//
			16'h01d9: data = 8'b00000000;	//
			16'h01da: data = 8'b00000000;	//
			16'h01db: data = 8'b00000000;	//
			16'h01dc: data = 8'b00000000;	//
			16'h01dd: data = 8'b00000000;	//
			16'h01de: data = 8'b00000000;	//
			16'h01df: data = 8'b00000000;	//
			// code x001e (rs) record separator
			16'h01e0: data = 8'b00000000;	//
			16'h01e1: data = 8'b00000000;	//
			16'h01e2: data = 8'b00000000;	//
			16'h01e3: data = 8'b00000000;	//
			16'h01e4: data = 8'b00000000;	//
			16'h01e5: data = 8'b00000000;	//
			16'h01e6: data = 8'b00000000;	//
			16'h01e7: data = 8'b00000000;	//
			16'h01e8: data = 8'b00000000;	//
			16'h01e9: data = 8'b00000000;	//
			16'h01ea: data = 8'b00000000;	//
			16'h01eb: data = 8'b00000000;	//
			16'h01ec: data = 8'b00000000;	//
			16'h01ed: data = 8'b00000000;	//
			16'h01ee: data = 8'b00000000;	//
			16'h01ef: data = 8'b00000000;	//
			// code x001f (us) unit separator
			16'h01f0: data = 8'b00000000;	//
			16'h01f1: data = 8'b00000000;	//
			16'h01f2: data = 8'b00000000;	//
			16'h01f3: data = 8'b00000000;	//
			16'h01f4: data = 8'b00000000;	//
			16'h01f5: data = 8'b00000000;	//
			16'h01f6: data = 8'b00000000;	//
			16'h01f7: data = 8'b00000000;	//
			16'h01f8: data = 8'b00000000;	//
			16'h01f9: data = 8'b00000000;	//
			16'h01fa: data = 8'b00000000;	//
			16'h01fb: data = 8'b00000000;	//
			16'h01fc: data = 8'b00000000;	//
			16'h01fd: data = 8'b00000000;	//
			16'h01fe: data = 8'b00000000;	//
			16'h01ff: data = 8'b00000000;	//		
		
			// Begin printable ASCII characters (20 -7e)
			// code x0020 ( ) -space-
			16'h0200: data = 8'b00000000;	//
			16'h0201: data = 8'b00000000;	//
			16'h0202: data = 8'b00000000;	//
			16'h0203: data = 8'b00000000;	//
			16'h0204: data = 8'b00000000;	//
			16'h0205: data = 8'b00000000;	//
			16'h0206: data = 8'b00000000;	//
			16'h0207: data = 8'b00000000;	//
			16'h0208: data = 8'b00000000;	//
			16'h0209: data = 8'b00000000;	//
			16'h020a: data = 8'b00000000;	//
			16'h020b: data = 8'b00000000;	//
			16'h020c: data = 8'b00000000;	//
			16'h020d: data = 8'b00000000;	//
			16'h020e: data = 8'b00000000;	//
			16'h020f: data = 8'b00000000;	//
			// code x0021 (!)
			16'h0210: data = 8'b00000000;	//
			16'h0211: data = 8'b00000000;	//
			16'h0212: data = 8'b00000000;	//
			16'h0213: data = 8'b00011000;	//   **
			16'h0214: data = 8'b00011000;	//   **
			16'h0215: data = 8'b00011000;	//   **
			16'h0216: data = 8'b00011000;	//   **
			16'h0217: data = 8'b00011000;	//   **
			16'h0218: data = 8'b00011000;	//   **
			16'h0219: data = 8'b00000000;	//
			16'h021a: data = 8'b00011000;	//   **
			16'h021b: data = 8'b00011000;	//   **
			16'h021c: data = 8'b00000000;	//
			16'h021d: data = 8'b00000000;	//
			16'h021e: data = 8'b00000000;	//
			16'h021f: data = 8'b00000000;	//
			// code x0022 (")
			16'h0220: data = 8'b00000000;	//
			16'h0221: data = 8'b00000000;	//
			16'h0222: data = 8'b00000000;	//
			16'h0223: data = 8'b00000000;	//
			16'h0224: data = 8'b00000000;	//
			16'h0225: data = 8'b00000000;	//
			16'h0226: data = 8'b00000000;	//
			16'h0227: data = 8'b00000000;	//
			16'h0228: data = 8'b00000000;	//
			16'h0229: data = 8'b00000000;	//
			16'h022a: data = 8'b00000000;	//
			16'h022b: data = 8'b00000000;	//
			16'h022c: data = 8'b00000000;	//
			16'h022d: data = 8'b00000000;	//
			16'h022e: data = 8'b00000000;	//
			16'h022f: data = 8'b00000000;	//
			// code x0023 (#)
			16'h0230: data = 8'b00000000;	//
			16'h0231: data = 8'b00000000;	//
			16'h0232: data = 8'b00000000;	//
			16'h0233: data = 8'b00000000;	//
			16'h0234: data = 8'b00000000;	//
			16'h0235: data = 8'b00000000;	//
			16'h0236: data = 8'b00000000;	//
			16'h0237: data = 8'b00000000;	//
			16'h0238: data = 8'b00000000;	//
			16'h0239: data = 8'b00000000;	//
			16'h023a: data = 8'b00000000;	//
			16'h023b: data = 8'b00000000;	//
			16'h023c: data = 8'b00000000;	//
			16'h023d: data = 8'b00000000;	//
			16'h023e: data = 8'b00000000;	//
			16'h023f: data = 8'b00000000;	//
			// code x0024 ($)
			16'h0240: data = 8'b00000000;	//
			16'h0241: data = 8'b00000000;	//
			16'h0242: data = 8'b00000000;	//
			16'h0243: data = 8'b00000000;	//
			16'h0244: data = 8'b00000000;	//
			16'h0245: data = 8'b00000000;	//
			16'h0246: data = 8'b00000000;	//
			16'h0247: data = 8'b00000000;	//
			16'h0248: data = 8'b00000000;	//
			16'h0249: data = 8'b00000000;	//
			16'h024a: data = 8'b00000000;	//
			16'h024b: data = 8'b00000000;	//
			16'h024c: data = 8'b00000000;	//
			16'h024d: data = 8'b00000000;	//
			16'h024e: data = 8'b00000000;	//
			16'h024f: data = 8'b00000000;	//
			// code x0025 (%)
			16'h0250: data = 8'b00000000;	//
			16'h0251: data = 8'b00000000;	//
			16'h0252: data = 8'b00000000;	//
			16'h0253: data = 8'b00000000;	//
			16'h0254: data = 8'b00000000;	//
			16'h0255: data = 8'b00000000;	//
			16'h0256: data = 8'b00000000;	//
			16'h0257: data = 8'b00000000;	//
			16'h0258: data = 8'b00000000;	//
			16'h0259: data = 8'b00000000;	//
			16'h025a: data = 8'b00000000;	//
			16'h025b: data = 8'b00000000;	//
			16'h025c: data = 8'b00000000;	//
			16'h025d: data = 8'b00000000;	//
			16'h025e: data = 8'b00000000;	//
			16'h025f: data = 8'b00000000;	//
			// code x0026 (&)
			16'h0260: data = 8'b00000000;	//
			16'h0261: data = 8'b00000000;	//
			16'h0262: data = 8'b00000000;	//
			16'h0263: data = 8'b00000000;	//
			16'h0264: data = 8'b00000000;	//
			16'h0265: data = 8'b00000000;	//
			16'h0266: data = 8'b00000000;	//
			16'h0267: data = 8'b00000000;	//
			16'h0268: data = 8'b00000000;	//
			16'h0269: data = 8'b00000000;	//
			16'h026a: data = 8'b00000000;	//
			16'h026b: data = 8'b00000000;	//
			16'h026c: data = 8'b00000000;	//
			16'h026d: data = 8'b00000000;	//
			16'h026e: data = 8'b00000000;	//
			16'h026f: data = 8'b00000000;	//
			// code x0027 (')
			16'h0270: data = 8'b00000000;	//
			16'h0271: data = 8'b00000000;	//
			16'h0272: data = 8'b00000000;	//
			16'h0273: data = 8'b00000000;	//
			16'h0274: data = 8'b00000000;	//
			16'h0275: data = 8'b00000000;	//
			16'h0276: data = 8'b00000000;	//
			16'h0277: data = 8'b00000000;	//
			16'h0278: data = 8'b00000000;	//
			16'h0279: data = 8'b00000000;	//
			16'h027a: data = 8'b00000000;	//
			16'h027b: data = 8'b00000000;	//
			16'h027c: data = 8'b00000000;	//
			16'h027d: data = 8'b00000000;	//
			16'h027e: data = 8'b00000000;	//
			16'h027f: data = 8'b00000000;	//
			// code x0028 (()
			16'h0280: data = 8'b00000000;	//
			16'h0281: data = 8'b00000000;	//
			16'h0282: data = 8'b00000000;	//
			16'h0283: data = 8'b00000000;	//
			16'h0284: data = 8'b00000000;	//
			16'h0285: data = 8'b00000000;	//
			16'h0286: data = 8'b00000000;	//
			16'h0287: data = 8'b00000000;	//
			16'h0288: data = 8'b00000000;	//
			16'h0289: data = 8'b00000000;	//
			16'h028a: data = 8'b00000000;	//
			16'h028b: data = 8'b00000000;	//
			16'h028c: data = 8'b00000000;	//
			16'h028d: data = 8'b00000000;	//
			16'h028e: data = 8'b00000000;	//
			16'h028f: data = 8'b00000000;	//
			// code x0029 ())
			16'h0290: data = 8'b00000000;	//
			16'h0291: data = 8'b00000000;	//
			16'h0292: data = 8'b00000000;	//
			16'h0293: data = 8'b00000000;	//
			16'h0294: data = 8'b00000000;	//
			16'h0295: data = 8'b00000000;	//
			16'h0296: data = 8'b00000000;	//
			16'h0297: data = 8'b00000000;	//
			16'h0298: data = 8'b00000000;	//
			16'h0299: data = 8'b00000000;	//
			16'h029a: data = 8'b00000000;	//
			16'h029b: data = 8'b00000000;	//
			16'h029c: data = 8'b00000000;	//
			16'h029d: data = 8'b00000000;	//
			16'h029e: data = 8'b00000000;	//
			16'h029f: data = 8'b00000000;	//
			// code x002a (*)
			16'h02a0: data = 8'b00000000;	//
			16'h02a1: data = 8'b00000000;	//
			16'h02a2: data = 8'b00000000;	//
			16'h02a3: data = 8'b00000000;	//
			16'h02a4: data = 8'b00000000;	//
			16'h02a5: data = 8'b00000000;	//
			16'h02a6: data = 8'b00000000;	//
			16'h02a7: data = 8'b00000000;	//
			16'h02a8: data = 8'b00000000;	//
			16'h02a9: data = 8'b00000000;	//
			16'h02aa: data = 8'b00000000;	//
			16'h02ab: data = 8'b00000000;	//
			16'h02ac: data = 8'b00000000;	//
			16'h02ad: data = 8'b00000000;	//
			16'h02ae: data = 8'b00000000;	//
			16'h02af: data = 8'b00000000;	//
			// code x002b (+)
			16'h02b0: data = 8'b00000000;	//
			16'h02b1: data = 8'b00000000;	//
			16'h02b2: data = 8'b00000000;	//
			16'h02b3: data = 8'b00010000;	//   *
			16'h02b4: data = 8'b00010000;	//   *
			16'h02b5: data = 8'b00010000;	//   *
			16'h02b6: data = 8'b11111110;	//*******
			16'h02b7: data = 8'b00010000;	//   *
			16'h02b8: data = 8'b00010000;	//   *
			16'h02b9: data = 8'b00010000;	//   *
			16'h02ba: data = 8'b00000000;	//
			16'h02bb: data = 8'b00000000;	//
			16'h02bc: data = 8'b00000000;	//
			16'h02bd: data = 8'b00000000;	//
			16'h02be: data = 8'b00000000;	//
			16'h02bf: data = 8'b00000000;	//
			// code x002c (,)
			16'h02c0: data = 8'b00000000;	//
			16'h02c1: data = 8'b00000000;	//
			16'h02c2: data = 8'b00000000;	//
			16'h02c3: data = 8'b00000000;	//
			16'h02c4: data = 8'b00000000;	//
			16'h02c5: data = 8'b00000000;	//
			16'h02c6: data = 8'b00000000;	//
			16'h02c7: data = 8'b00000000;	//
			16'h02c8: data = 8'b00000000;	//
			16'h02c9: data = 8'b00000000;	//
			16'h02ca: data = 8'b00000000;	//
			16'h02cb: data = 8'b00000000;	//
			16'h02cc: data = 8'b00000000;	//
			16'h02cd: data = 8'b00000000;	//
			16'h02ce: data = 8'b00000000;	//
			16'h02cf: data = 8'b00000000;	//
			// code x002d (-)
			16'h02d0: data = 8'b00000000;	//
			16'h02d1: data = 8'b00000000;	//
			16'h02d2: data = 8'b00000000;	//
			16'h02d3: data = 8'b00000000;	//
			16'h02d4: data = 8'b00000000;	//
			16'h02d5: data = 8'b00000000;	//
			16'h02d6: data = 8'b01111110;	// ******
			16'h02d7: data = 8'b00000000;	//
			16'h02d8: data = 8'b00000000;	//
			16'h02d9: data = 8'b00000000;	//
			16'h02da: data = 8'b00000000;	//
			16'h02db: data = 8'b00000000;	//
			16'h02dc: data = 8'b00000000;	//
			16'h02dd: data = 8'b00000000;	//
			16'h02de: data = 8'b00000000;	//
			16'h02df: data = 8'b00000000;	//
			// code x002e (.)
			16'h02e0: data = 8'b00000000;	//
			16'h02e1: data = 8'b00000000;	//
			16'h02e2: data = 8'b00000000;	//
			16'h02e3: data = 8'b00000000;	//
			16'h02e4: data = 8'b00000000;	//
			16'h02e5: data = 8'b00000000;	//
			16'h02e6: data = 8'b00000000;	//
			16'h02e7: data = 8'b00000000;	//
			16'h02e8: data = 8'b00000000;	//
			16'h02e9: data = 8'b00000000;	//
			16'h02ea: data = 8'b00011000;	//   **
			16'h02eb: data = 8'b00011000;	//   **
			16'h02ec: data = 8'b00000000;	//
			16'h02ed: data = 8'b00000000;	//
			16'h02ee: data = 8'b00000000;	//
			16'h02ef: data = 8'b00000000;	//
			// code x002f (/)
			16'h02f0: data = 8'b00000000;	//
			16'h02f1: data = 8'b00000000;	//
			16'h02f2: data = 8'b00000000;	//
			16'h02f3: data = 8'b00000000;	//
			16'h02f4: data = 8'b00000000;	//
			16'h02f5: data = 8'b00000000;	//
			16'h02f6: data = 8'b00000000;	//
			16'h02f7: data = 8'b00000000;	//
			16'h02f8: data = 8'b00000000;	//
			16'h02f9: data = 8'b00000000;	//
			16'h02fa: data = 8'b00000000;	//
			16'h02fb: data = 8'b00000000;	//
			16'h02fc: data = 8'b00000000;	//
			16'h02fd: data = 8'b00000000;	//
			16'h02fe: data = 8'b00000000;	//
			16'h02ff: data = 8'b00000000;	//
			// code x0030 (0)
			16'h0300: data = 8'b00000000;	//
			16'h0301: data = 8'b00000000;	//
			16'h0302: data = 8'b00111000;	//  ***  
			16'h0303: data = 8'b01101100;	// ** **
			16'h0304: data = 8'b11000110;	//**   **
			16'h0305: data = 8'b11000110;	//**   **
			16'h0306: data = 8'b11000110;	//**   **
			16'h0307: data = 8'b11000110;	//**   **
			16'h0308: data = 8'b11000110;	//**   **
			16'h0309: data = 8'b11000110;	//**   **
			16'h030a: data = 8'b01101100;	// ** **
			16'h030b: data = 8'b00111000;	//  ***
			16'h030c: data = 8'b00000000;	//
			16'h030d: data = 8'b00000000;	//
			16'h030e: data = 8'b00000000;	//
			16'h030f: data = 8'b00000000;	//
			// code x0031 (1)
			16'h0310: data = 8'b00000000;	//
			16'h0311: data = 8'b00000000;	//
			16'h0312: data = 8'b00011000;	//   **  
			16'h0313: data = 8'b00111000;	//  ***
			16'h0314: data = 8'b01111000;	// ****
			16'h0315: data = 8'b00011000;	//   **
			16'h0316: data = 8'b00011000;	//   **
			16'h0317: data = 8'b00011000;	//   **
			16'h0318: data = 8'b00011000;	//   **
			16'h0319: data = 8'b00011000;	//   **
			16'h031a: data = 8'b01111110;	// ******
			16'h031b: data = 8'b01111110;	// ******
			16'h031c: data = 8'b00000000;	//
			16'h031d: data = 8'b00000000;	//
			16'h031e: data = 8'b00000000;	//
			16'h031f: data = 8'b00000000;	//
			// code x0032 (2)
			16'h0320: data = 8'b00000000;	//
			16'h0321: data = 8'b00000000;	//
			16'h0322: data = 8'b11111110;	//*******  
			16'h0323: data = 8'b11111110;	//*******
			16'h0324: data = 8'b00000110;	//     **
			16'h0325: data = 8'b00000110;	//     **
			16'h0326: data = 8'b11111110;	//*******
			16'h0327: data = 8'b11111110;	//*******
			16'h0328: data = 8'b11000000;	//**
			16'h0329: data = 8'b11000000;	//**
			16'h032a: data = 8'b11111110;	//*******
			16'h032b: data = 8'b11111110;	//*******
			16'h032c: data = 8'b00000000;	//
			16'h032d: data = 8'b00000000;	//
			16'h032e: data = 8'b00000000;	//
			16'h032f: data = 8'b00000000;	//
			// code x0033 (3)
			16'h0330: data = 8'b00000000;	//
			16'h0331: data = 8'b00000000;	//
			16'h0332: data = 8'b11111110;	//*******  
			16'h0333: data = 8'b11111110;	//*******
			16'h0334: data = 8'b00000110;	//     **
			16'h0335: data = 8'b00000110;	//     **
			16'h0336: data = 8'b00111110;	//  *****
			16'h0337: data = 8'b00111110;	//  *****
			16'h0338: data = 8'b00000110;	//     **
			16'h0339: data = 8'b00000110;	//     **
			16'h033a: data = 8'b11111110;	//*******
			16'h033b: data = 8'b11111110;	//*******
			16'h033c: data = 8'b00000000;	//
			16'h033d: data = 8'b00000000;	//
			16'h033e: data = 8'b00000000;	//
			16'h033f: data = 8'b00000000;	//
			// code x0034 (4)
			16'h0340: data = 8'b00000000;	//
			16'h0341: data = 8'b00000000;	//
			16'h0342: data = 8'b11000110;	//**   **  
			16'h0343: data = 8'b11000110;	//**   **
			16'h0344: data = 8'b11000110;	//**   **
			16'h0345: data = 8'b11000110;	//**   **
			16'h0346: data = 8'b11111110;	//*******
			16'h0347: data = 8'b11111110;	//*******
			16'h0348: data = 8'b00000110;	//     **
			16'h0349: data = 8'b00000110;	//     **
			16'h034a: data = 8'b00000110;	//     **
			16'h034b: data = 8'b00000110;	//     **
			16'h034c: data = 8'b00000000;	//
			16'h034d: data = 8'b00000000;	//
			16'h034e: data = 8'b00000000;	//
			16'h034f: data = 8'b00000000;	//
			// code x0035 (5)
			16'h0350: data = 8'b00000000;	//
			16'h0351: data = 8'b00000000;	//
			16'h0352: data = 8'b11111110;	//*******  
			16'h0353: data = 8'b11111110;	//*******
			16'h0354: data = 8'b11000000;	//**
			16'h0355: data = 8'b11000000;	//**
			16'h0356: data = 8'b11111110;	//*******
			16'h0357: data = 8'b11111110;	//*******
			16'h0358: data = 8'b00000110;	//     **
			16'h0359: data = 8'b00000110;	//     **
			16'h035a: data = 8'b11111110;	//*******
			16'h035b: data = 8'b11111110;	//*******
			16'h035c: data = 8'b00000000;	//
			16'h035d: data = 8'b00000000;	//
			16'h035e: data = 8'b00000000;	//
			16'h035f: data = 8'b00000000;	//
			// code x0036 (6)
			16'h0360: data = 8'b00000000;	//
			16'h0361: data = 8'b00000000;	//
			16'h0362: data = 8'b11111110;	//*******  
			16'h0363: data = 8'b11111110;	//*******
			16'h0364: data = 8'b11000000;	//**
			16'h0365: data = 8'b11000000;	//**
			16'h0366: data = 8'b11111110;	//*******
			16'h0367: data = 8'b11111110;	//*******
			16'h0368: data = 8'b11000110;	//**   **
			16'h0369: data = 8'b11000110;	//**   **
			16'h036a: data = 8'b11111110;	//*******
			16'h036b: data = 8'b11111110;	//*******
			16'h036c: data = 8'b00000000;	//
			16'h036d: data = 8'b00000000;	//
			16'h036e: data = 8'b00000000;	//
			16'h036f: data = 8'b00000000;	//
			// code x0037 (7)
			16'h0370: data = 8'b00000000;	//
			16'h0371: data = 8'b00000000;	//
			16'h0372: data = 8'b11111110;	//*******  
			16'h0373: data = 8'b11111110;	//*******
			16'h0374: data = 8'b00000110;	//     **
			16'h0375: data = 8'b00000110;	//     **
			16'h0376: data = 8'b00000110;	//     **
			16'h0377: data = 8'b00000110;	//     **
			16'h0378: data = 8'b00000110;	//     **
			16'h0379: data = 8'b00000110;	//     **
			16'h037a: data = 8'b00000110;	//     **
			16'h037b: data = 8'b00000110;	//     **
			16'h037c: data = 8'b00000000;	//
			16'h037d: data = 8'b00000000;	//
			16'h037e: data = 8'b00000000;	//
			16'h037f: data = 8'b00000000;	//
			// code x0038 (8)
			16'h0380: data = 8'b00000000;	//
			16'h0381: data = 8'b00000000;	//
			16'h0382: data = 8'b11111110;	//*******  
			16'h0383: data = 8'b11111110;	//*******
			16'h0384: data = 8'b11000110;	//**   **
			16'h0385: data = 8'b11000110;	//**   **
			16'h0386: data = 8'b11111110;	//*******
			16'h0387: data = 8'b11111110;	//*******
			16'h0388: data = 8'b11000110;	//**   **
			16'h0389: data = 8'b11000110;	//**   **
			16'h038a: data = 8'b11111110;	//*******
			16'h038b: data = 8'b11111110;	//*******
			16'h038c: data = 8'b00000000;	//
			16'h038d: data = 8'b00000000;	//
			16'h038e: data = 8'b00000000;	//
			16'h038f: data = 8'b00000000;	//
			// code x0039 (9)
			16'h0390: data = 8'b00000000;	//
			16'h0391: data = 8'b00000000;	//
			16'h0392: data = 8'b11111110;	//*******  
			16'h0393: data = 8'b11111110;	//*******
			16'h0394: data = 8'b11000110;	//**   **
			16'h0395: data = 8'b11000110;	//**   **
			16'h0396: data = 8'b11111110;	//*******
			16'h0397: data = 8'b11111110;	//*******
			16'h0398: data = 8'b00000110;	//     **
			16'h0399: data = 8'b00000110;	//     **
			16'h039a: data = 8'b11111110;	//*******
			16'h039b: data = 8'b11111110;	//*******
			16'h039c: data = 8'b00000000;	//
			16'h039d: data = 8'b00000000;	//
			16'h039e: data = 8'b00000000;	//
			16'h039f: data = 8'b00000000;	//
			// code x003a (:)
			16'h03a0: data = 8'b00000000;	//
			16'h03a1: data = 8'b00000000;	//
			16'h03a2: data = 8'b00000000;	//
			16'h03a3: data = 8'b00000000;	//
			16'h03a4: data = 8'b00011000;	//   **
			16'h03a5: data = 8'b00011000;	//   **
			16'h03a6: data = 8'b00000000;	//
			16'h03a7: data = 8'b00000000;	//
			16'h03a8: data = 8'b00011000;	//   **
			16'h03a9: data = 8'b00011000;	//   **
			16'h03aa: data = 8'b00000000;	//   
			16'h03ab: data = 8'b00000000;	//   
			16'h03ac: data = 8'b00000000;	//
			16'h03ad: data = 8'b00000000;	//
			16'h03ae: data = 8'b00000000;	//
			16'h03af: data = 8'b00000000;	//
			// code x003b (;)
			16'h03b0: data = 8'b00000000;	//
			16'h03b1: data = 8'b00000000;	//
			16'h03b2: data = 8'b00000000;	//
			16'h03b3: data = 8'b00000000;	//
			16'h03b4: data = 8'b00000000;	//
			16'h03b5: data = 8'b00000000;	//
			16'h03b6: data = 8'b00000000;	//
			16'h03b7: data = 8'b00000000;	//
			16'h03b8: data = 8'b00000000;	//
			16'h03b9: data = 8'b00000000;	//
			16'h03ba: data = 8'b00000000;	//
			16'h03bb: data = 8'b00000000;	//
			16'h03bc: data = 8'b00000000;	//
			16'h03bd: data = 8'b00000000;	//
			16'h03be: data = 8'b00000000;	//
			16'h03bf: data = 8'b00000000;	//
			// code x003c (<)
			16'h03c0: data = 8'b00000000;	//
			16'h03c1: data = 8'b00000000;	//
			16'h03c2: data = 8'b00000000;	//
			16'h03c3: data = 8'b00000000;	//
			16'h03c4: data = 8'b00000000;	//
			16'h03c5: data = 8'b00000000;	//
			16'h03c6: data = 8'b00000000;	//
			16'h03c7: data = 8'b00000000;	//
			16'h03c8: data = 8'b00000000;	//
			16'h03c9: data = 8'b00000000;	//
			16'h03ca: data = 8'b00000000;	//
			16'h03cb: data = 8'b00000000;	//
			16'h03cc: data = 8'b00000000;	//
			16'h03cd: data = 8'b00000000;	//
			16'h03ce: data = 8'b00000000;	//
			16'h03cf: data = 8'b00000000;	//
			// code x003d (=)
			16'h03d0: data = 8'b00000000;	//
			16'h03d1: data = 8'b00000000;	//
			16'h03d2: data = 8'b00000000;	//
			16'h03d3: data = 8'b00000000;	//
			16'h03d4: data = 8'b00000000;	//
			16'h03d5: data = 8'b00000000;	//
			16'h03d6: data = 8'b01111110;	// ******
			16'h03d7: data = 8'b00000000;	// 
			16'h03d8: data = 8'b01111110;	// ******
			16'h03d9: data = 8'b00000000;	//
			16'h03da: data = 8'b00000000;	//
			16'h03db: data = 8'b00000000;	//
			16'h03dc: data = 8'b00000000;	//
			16'h03dd: data = 8'b00000000;	//
			16'h03de: data = 8'b00000000;	//
			16'h03df: data = 8'b00000000;	//
			// code x003e (>)
			16'h03e0: data = 8'b00000000;	//
			16'h03e1: data = 8'b00000000;	//
			16'h03e2: data = 8'b00000000;	//
			16'h03e3: data = 8'b00000000;	//
			16'h03e4: data = 8'b00000000;	//
			16'h03e5: data = 8'b00000000;	//
			16'h03e6: data = 8'b00000000;	//
			16'h03e7: data = 8'b00000000;	//
			16'h03e8: data = 8'b00000000;	//
			16'h03e9: data = 8'b00000000;	//
			16'h03ea: data = 8'b00000000;	//
			16'h03eb: data = 8'b00000000;	//
			16'h03ec: data = 8'b00000000;	//
			16'h03ed: data = 8'b00000000;	//
			16'h03ee: data = 8'b00000000;	//
			16'h03ef: data = 8'b00000000;	//
			// code x003f (?)
			16'h03f0: data = 8'b00000000;	//
			16'h03f1: data = 8'b00000000;	//
			16'h03f2: data = 8'b00000000;	//
			16'h03f3: data = 8'b00000000;	//
			16'h03f4: data = 8'b00000000;	//
			16'h03f5: data = 8'b00000000;	//
			16'h03f6: data = 8'b00000000;	//
			16'h03f7: data = 8'b00000000;	//
			16'h03f8: data = 8'b00000000;	//
			16'h03f9: data = 8'b00000000;	//
			16'h03fa: data = 8'b00000000;	//
			16'h03fb: data = 8'b00000000;	//
			16'h03fc: data = 8'b00000000;	//
			16'h03fd: data = 8'b00000000;	//
			16'h03fe: data = 8'b00000000;	//
			16'h03ff: data = 8'b00000000;	//
			// code x0040 (@)
			16'h0400: data = 8'b00000000;	//
			16'h0401: data = 8'b00000000;	//
			16'h0402: data = 8'b00000000;	//
			16'h0403: data = 8'b00000000;	//
			16'h0404: data = 8'b00000000;	//
			16'h0405: data = 8'b00000000;	//
			16'h0406: data = 8'b00000000;	//
			16'h0407: data = 8'b00000000;	//
			16'h0408: data = 8'b00000000;	//
			16'h0409: data = 8'b00000000;	//
			16'h040a: data = 8'b00000000;	//
			16'h040b: data = 8'b00000000;	//
			16'h040c: data = 8'b00000000;	//
			16'h040d: data = 8'b00000000;	//
			16'h040e: data = 8'b00000000;	//
			16'h040f: data = 8'b00000000;	//		
			// code x0041 (A)
			16'h0410: data = 8'b00000000;	//
			16'h0411: data = 8'b00000000;	//
			16'h0412: data = 8'b00010000;	//   *
			16'h0413: data = 8'b00111000;	//  ***
			16'h0414: data = 8'b01101100;	// ** **   
			16'h0415: data = 8'b11000110;	//**   **   
			16'h0416: data = 8'b11000110;	//**   **
			16'h0417: data = 8'b11111110;	//*******
			16'h0418: data = 8'b11111110;	//*******
			16'h0419: data = 8'b11000110;	//**   **
			16'h041a: data = 8'b11000110;	//**   **
			16'h041b: data = 8'b11000110;	//**   **
			16'h041c: data = 8'b00000000;	//
			16'h041d: data = 8'b00000000;	//
			16'h041e: data = 8'b00000000;	//
			16'h041f: data = 8'b00000000;	//
			// code x0042 (B)
			16'h0420: data = 8'b00000000;	//
			16'h0421: data = 8'b00000000;	//
			16'h0422: data = 8'b11111100;	//******
			16'h0423: data = 8'b11111110;	//*******
			16'h0424: data = 8'b11000110;	//**   **
			16'h0425: data = 8'b11000110;	//**   **   
			16'h0426: data = 8'b11111100;	//******
			16'h0427: data = 8'b11111100;	//******
			16'h0428: data = 8'b11000110;	//**   **
			16'h0429: data = 8'b11000110;	//**   **
			16'h042a: data = 8'b11111110;	//*******
			16'h042b: data = 8'b11111100;	//******
			16'h042c: data = 8'b00000000;	//
			16'h042d: data = 8'b00000000;	//
			16'h042e: data = 8'b00000000;	//
			16'h042f: data = 8'b00000000;	//
			// code x0043 (C)
			16'h0430: data = 8'b00000000;	//
			16'h0431: data = 8'b00000000;	//
			16'h0432: data = 8'b01111100;	// *****
			16'h0433: data = 8'b11111110;	//*******
			16'h0434: data = 8'b11000000;	//**
			16'h0435: data = 8'b11000000;	//**   
			16'h0436: data = 8'b11000000;	//**
			16'h0437: data = 8'b11000000;	//**
			16'h0438: data = 8'b11000000;	//** 
			16'h0439: data = 8'b11000000;	//** 
			16'h043a: data = 8'b11111110;	//*******
			16'h043b: data = 8'b01111100;	// *****
			16'h043c: data = 8'b00000000;	//
			16'h043d: data = 8'b00000000;	//
			16'h043e: data = 8'b00000000;	//
			16'h043f: data = 8'b00000000;	//
			// code x0044 (D)
			16'h0440: data = 8'b00000000;	//
			16'h0441: data = 8'b00000000;	//
			16'h0442: data = 8'b11111100;	//******
			16'h0443: data = 8'b11111110;	//*******
			16'h0444: data = 8'b11000110;	//**   **
			16'h0445: data = 8'b11000110;	//**   **   
			16'h0446: data = 8'b11000110;	//**   **
			16'h0447: data = 8'b11000110;	//**   **
			16'h0448: data = 8'b11000110;	//**   ** 
			16'h0449: data = 8'b11000110;	//**   ** 
			16'h044a: data = 8'b11111110;	//*******
			16'h044b: data = 8'b11111100;	//******
			16'h044c: data = 8'b00000000;	//
			16'h044d: data = 8'b00000000;	//
			16'h044e: data = 8'b00000000;	//
			16'h044f: data = 8'b00000000;	//
			// code x0045 (E)
			16'h0450: data = 8'b00000000;	//
			16'h0451: data = 8'b00000000;	//
			16'h0452: data = 8'b11111110;	//*******
			16'h0453: data = 8'b11111110;	//*******
			16'h0454: data = 8'b11000000;	//**
			16'h0455: data = 8'b11000000;	//**   
			16'h0456: data = 8'b11111100;	//******
			16'h0457: data = 8'b11111100;	//******
			16'h0458: data = 8'b11000000;	//** 
			16'h0459: data = 8'b11000000;	//** 
			16'h045a: data = 8'b11111110;	//*******
			16'h045b: data = 8'b11111110;	//*******
			16'h045c: data = 8'b00000000;	//
			16'h045d: data = 8'b00000000;	//
			16'h045e: data = 8'b00000000;	//
			16'h045f: data = 8'b00000000;	//
			// code x0046 (F)
			16'h0460: data = 8'b00000000;	//
			16'h0461: data = 8'b00000000;	//
			16'h0462: data = 8'b11111110;	//*******
			16'h0463: data = 8'b11111110;	//*******
			16'h0464: data = 8'b11000000;	//**
			16'h0465: data = 8'b11000000;	//**   
			16'h0466: data = 8'b11111100;	//******
			16'h0467: data = 8'b11111100;	//******
			16'h0468: data = 8'b11000000;	//** 
			16'h0469: data = 8'b11000000;	//** 
			16'h046a: data = 8'b11000000;	//**
			16'h046b: data = 8'b11000000;	//**
			16'h046c: data = 8'b00000000;	//
			16'h046d: data = 8'b00000000;	//
			16'h046e: data = 8'b00000000;	//
			16'h046f: data = 8'b00000000;	//
			// code x0047 (G)
			16'h0470: data = 8'b00000000;	//
			16'h0471: data = 8'b00000000;	//
			16'h0472: data = 8'b01111100;	// *****
			16'h0473: data = 8'b11111110;	//*******
			16'h0474: data = 8'b11000000;	//**
			16'h0475: data = 8'b11000000;	//**   
			16'h0476: data = 8'b11111110;	//*******
			16'h0477: data = 8'b11111110;	//*******
			16'h0478: data = 8'b11000110;	//**   **
			16'h0479: data = 8'b11000110;	//**   **
			16'h047a: data = 8'b11111110;	//*******
			16'h047b: data = 8'b01110110;	// *** **
			16'h047c: data = 8'b00000000;	//
			16'h047d: data = 8'b00000000;	//
			16'h047e: data = 8'b00000000;	//
			16'h047f: data = 8'b00000000;	//
			// code x0048 (H)
			16'h0480: data = 8'b00000000;	//
			16'h0481: data = 8'b00000000;	//
			16'h0482: data = 8'b11000110;	//**   **
			16'h0483: data = 8'b11000110;	//**   **
			16'h0484: data = 8'b11000110;	//**   **
			16'h0485: data = 8'b11000110;	//**   **
			16'h0486: data = 8'b11111110;	//*******
			16'h0487: data = 8'b11111110;	//*******
			16'h0488: data = 8'b11000110;	//**   **
			16'h0489: data = 8'b11000110;	//**   **
			16'h048a: data = 8'b11000110;	//**   **
			16'h048b: data = 8'b11000110;	//**   **
			16'h048c: data = 8'b00000000;	//
			16'h048d: data = 8'b00000000;	//
			16'h048e: data = 8'b00000000;	//
			16'h048f: data = 8'b00000000;	//
			// code x0049 (I)
			16'h0490: data = 8'b00000000;	//
			16'h0491: data = 8'b00000000;	//
			16'h0492: data = 8'b11111110;	//*******
			16'h0493: data = 8'b11111110;	//*******
			16'h0494: data = 8'b00110000;	//  **
			16'h0495: data = 8'b00110000;	//  **
			16'h0496: data = 8'b00110000;	//  **
			16'h0497: data = 8'b00110000;	//  **
			16'h0498: data = 8'b00110000;	//  **
			16'h0499: data = 8'b00110000;	//  **
			16'h049a: data = 8'b11111110;	//*******
			16'h049b: data = 8'b11111110;	//*******
			16'h049c: data = 8'b00000000;	//
			16'h049d: data = 8'b00000000;	//
			16'h049e: data = 8'b00000000;	//
			16'h049f: data = 8'b00000000;	//
			// code x004a (J)
			16'h04a0: data = 8'b00000000;	//
			16'h04a1: data = 8'b00000000;	//
			16'h04a2: data = 8'b11111110;	//*******
			16'h04a3: data = 8'b11111110;	//*******
			16'h04a4: data = 8'b00011000;	//   **
			16'h04a5: data = 8'b00011000;	//   **
			16'h04a6: data = 8'b00011000;	//   **
			16'h04a7: data = 8'b00011000;	//   **
			16'h04a8: data = 8'b00011000;	//   **
			16'h04a9: data = 8'b00011000;	//   **
			16'h04aa: data = 8'b11111000;	//*****
			16'h04ab: data = 8'b01111000;	// ****
			16'h04ac: data = 8'b00000000;	//
			16'h04ad: data = 8'b00000000;	//
			16'h04ae: data = 8'b00000000;	//
			16'h04af: data = 8'b00000000;	//
			// code x004b (K)
			16'h04b0: data = 8'b00000000;	//
			16'h04b1: data = 8'b00000000;	//
			16'h04b2: data = 8'b11000110;	//**   **
			16'h04b3: data = 8'b11001100;	//**  **
			16'h04b4: data = 8'b11011000;	//** **
			16'h04b5: data = 8'b11110000;	//****
			16'h04b6: data = 8'b11100000;	//***
			16'h04b7: data = 8'b11100000;	//***
			16'h04b8: data = 8'b11110000;	//****
			16'h04b9: data = 8'b11011000;	//** **
			16'h04ba: data = 8'b11001100;	//**  **
			16'h04bb: data = 8'b11000110;	//**   **
			16'h04bc: data = 8'b00000000;	//
			16'h04bd: data = 8'b00000000;	//
			16'h04be: data = 8'b00000000;	//
			16'h04bf: data = 8'b00000000;	//
			// code x004c (L)
			16'h04c0: data = 8'b00000000;	//
			16'h04c1: data = 8'b00000000;	//
			16'h04c2: data = 8'b11000000;	//**
			16'h04c3: data = 8'b11000000;	//**
			16'h04c4: data = 8'b11000000;	//**
			16'h04c5: data = 8'b11000000;	//**
			16'h04c6: data = 8'b11000000;	//**
			16'h04c7: data = 8'b11000000;	//**
			16'h04c8: data = 8'b11000000;	//**
			16'h04c9: data = 8'b11000000;	//**
			16'h04ca: data = 8'b11111110;	//*******
			16'h04cb: data = 8'b11111110;	//*******
			16'h04cc: data = 8'b00000000;	//
			16'h04cd: data = 8'b00000000;	//
			16'h04ce: data = 8'b00000000;	//
			16'h04cf: data = 8'b00000000;	//
			// code x004d (M)
			16'h04d0: data = 8'b00000000;	//
			16'h04d1: data = 8'b00000000;	//
			16'h04d2: data = 8'b11000110;	//**   **
			16'h04d3: data = 8'b11000110;	//**   **
			16'h04d4: data = 8'b11101110;	//*** ***
			16'h04d5: data = 8'b11111110;	//*******
			16'h04d6: data = 8'b11010110;	//** * **
			16'h04d7: data = 8'b11000110;	//**   **
			16'h04d8: data = 8'b11000110;	//**   **
			16'h04d9: data = 8'b11000110;	//**   **
			16'h04da: data = 8'b11000110;	//**   **
			16'h04db: data = 8'b11000110;	//**   **
			16'h04dc: data = 8'b00000000;	//
			16'h04dd: data = 8'b00000000;	//
			16'h04de: data = 8'b00000000;	//
			16'h04df: data = 8'b00000000;	//
			// code x004e (N)
			16'h04e0: data = 8'b00000000;	//
			16'h04e1: data = 8'b00000000;	//
			16'h04e2: data = 8'b11000110;	//**   **
			16'h04e3: data = 8'b11000110;	//**   **
			16'h04e4: data = 8'b11100110;	//***  **
			16'h04e5: data = 8'b11110110;	//**** **
			16'h04e6: data = 8'b11111110;	//*******
			16'h04e7: data = 8'b11011110;	//** ****
			16'h04e8: data = 8'b11001110;	//**  ***
			16'h04e9: data = 8'b11000110;	//**   **
			16'h04ea: data = 8'b11000110;	//**   **
			16'h04eb: data = 8'b11000110;	//**   **
			16'h04ec: data = 8'b00000000;	//
			16'h04ed: data = 8'b00000000;	//
			16'h04ee: data = 8'b00000000;	//
			16'h04ef: data = 8'b00000000;	//
			// code x004f (O)
			16'h04f0: data = 8'b00000000;	//
			16'h04f1: data = 8'b00000000;	//
			16'h04f2: data = 8'b01111100;	// *****
			16'h04f3: data = 8'b11111110;	//*******
			16'h04f4: data = 8'b11000110;	//**   **
			16'h04f5: data = 8'b11000110;	//**   **
			16'h04f6: data = 8'b11000110;	//**   **
			16'h04f7: data = 8'b11000110;	//**   **
			16'h04f8: data = 8'b11000110;	//**   **
			16'h04f9: data = 8'b11000110;	//**   **
			16'h04fa: data = 8'b11111110;	//*******
			16'h04fb: data = 8'b01111100;	// *****
			16'h04fc: data = 8'b00000000;	//
			16'h04fd: data = 8'b00000000;	//
			16'h04fe: data = 8'b00000000;	//
			16'h04ff: data = 8'b00000000;	//
			// code x0050 (P)
			16'h0500: data = 8'b00000000;	//
			16'h0501: data = 8'b00000000;	//
			16'h0502: data = 8'b11111100;	//******
			16'h0503: data = 8'b11111110;	//*******
			16'h0504: data = 8'b11000110;	//**   **
			16'h0505: data = 8'b11000110;	//**   **
			16'h0506: data = 8'b11111110;	//*******
			16'h0507: data = 8'b11111100;	//******   
			16'h0508: data = 8'b11000000;	//**   
			16'h0509: data = 8'b11000000;	//**   
			16'h050a: data = 8'b11000000;	//**
			16'h050b: data = 8'b11000000;	//**
			16'h050c: data = 8'b00000000;	//
			16'h050d: data = 8'b00000000;	//
			16'h050e: data = 8'b00000000;	//
			16'h050f: data = 8'b00000000;	//
			// code x0051 (Q)
			16'h0510: data = 8'b00000000;	//
			16'h0511: data = 8'b00000000;	//
			16'h0512: data = 8'b11111100;	// *****
			16'h0513: data = 8'b11111110;	//*******
			16'h0514: data = 8'b11000110;	//**   **
			16'h0515: data = 8'b11000110;	//**   **
			16'h0516: data = 8'b11000110;	//**   **
			16'h0517: data = 8'b11000110;	//**   **  
			16'h0518: data = 8'b11010110;	//** * **
			16'h0519: data = 8'b11111110;	//*******
			16'h051a: data = 8'b01101100;	// ** ** 
			16'h051b: data = 8'b00000110;	//     **
			16'h051c: data = 8'b00000000;	//
			16'h051d: data = 8'b00000000;	//
			16'h051e: data = 8'b00000000;	//
			16'h051f: data = 8'b00000000;	//
			// code x0052 (R)
			16'h0520: data = 8'b00000000;	//
			16'h0521: data = 8'b00000000;	//
			16'h0522: data = 8'b11111100;	//******
			16'h0523: data = 8'b11111110;	//*******
			16'h0524: data = 8'b11000110;	//**   **
			16'h0525: data = 8'b11000110;	//**   **
			16'h0526: data = 8'b11111110;	//*******
			16'h0527: data = 8'b11111100;	//******   
			16'h0528: data = 8'b11011000;	//** **  
			16'h0529: data = 8'b11001100;	//**  ** 
			16'h052a: data = 8'b11000110;	//**   **
			16'h052b: data = 8'b11000110;	//**   **
			16'h052c: data = 8'b00000000;	//
			16'h052d: data = 8'b00000000;	//
			16'h052e: data = 8'b00000000;	//
			16'h052f: data = 8'b00000000;	//
			// code x0053 (S)
			16'h0530: data = 8'b00000000;	//
			16'h0531: data = 8'b00000000;	//
			16'h0532: data = 8'b01111100;	// *****
			16'h0533: data = 8'b11111110;	//*******
			16'h0534: data = 8'b11000000;	//**   
			16'h0535: data = 8'b11000000;	//**   
			16'h0536: data = 8'b11111100;	//******
			16'h0537: data = 8'b01111110;	// ******   
			16'h0538: data = 8'b00000110;	//     **  
			16'h0539: data = 8'b00000110;	//     **
			16'h053a: data = 8'b11111110;	//*******  
			16'h053b: data = 8'b01111100;	// ***** 
			16'h053c: data = 8'b00000000;	//
			16'h053d: data = 8'b00000000;	//
			16'h053e: data = 8'b00000000;	//
			16'h053f: data = 8'b00000000;	//
			// code x0054 (T)
			16'h0540: data = 8'b00000000;	//
			16'h0541: data = 8'b00000000;	//
			16'h0542: data = 8'b11111110;	//*******
			16'h0543: data = 8'b11111110;	//*******
			16'h0544: data = 8'b00110000;	//  **
			16'h0545: data = 8'b00110000;	//  **
			16'h0546: data = 8'b00110000;	//  **
			16'h0547: data = 8'b00110000;	//  **   
			16'h0548: data = 8'b00110000;	//  **  
			16'h0549: data = 8'b00110000;	//  **
			16'h054a: data = 8'b00110000;	//  **  
			16'h054b: data = 8'b00110000;	//  **
			16'h054c: data = 8'b00000000;	//
			16'h054d: data = 8'b00000000;	//
			16'h054e: data = 8'b00000000;	//
			16'h054f: data = 8'b00000000;	//
			// code x0055 (U)
			16'h0550: data = 8'b00000000;	//
			16'h0551: data = 8'b00000000;	//
			16'h0552: data = 8'b11000110;	//**   **
			16'h0553: data = 8'b11000110;	//**   **
			16'h0554: data = 8'b11000110;	//**   **
			16'h0555: data = 8'b11000110;	//**   **
			16'h0556: data = 8'b11000110;	//**   **
			16'h0557: data = 8'b11000110;	//**   **
			16'h0558: data = 8'b11000110;	//**   **
			16'h0559: data = 8'b11000110;	//**   **
			16'h055a: data = 8'b11111110;	//*******
			16'h055b: data = 8'b01111100;	// *****
			16'h055c: data = 8'b00000000;	//
			16'h055d: data = 8'b00000000;	//
			16'h055e: data = 8'b00000000;	//
			16'h055f: data = 8'b00000000;	//
			// code x0056 (V)
			16'h0560: data = 8'b00000000;	//
			16'h0561: data = 8'b00000000;	//
			16'h0562: data = 8'b11000110;	//**   **
			16'h0563: data = 8'b11000110;	//**   **
			16'h0564: data = 8'b11000110;	//**   **
			16'h0565: data = 8'b11000110;	//**   **
			16'h0566: data = 8'b11000110;	//**   **
			16'h0567: data = 8'b11000110;	//**   **
			16'h0568: data = 8'b11000110;	//**   **
			16'h0569: data = 8'b01101100;	// ** **
			16'h056a: data = 8'b00111000;	//  ***  
			16'h056b: data = 8'b00010000;	//   * 
			16'h056c: data = 8'b00000000;	//
			16'h056d: data = 8'b00000000;	//
			16'h056e: data = 8'b00000000;	//
			16'h056f: data = 8'b00000000;	//
			// code x0057 (W)
			16'h0570: data = 8'b00000000;	//
			16'h0571: data = 8'b00000000;	//
			16'h0572: data = 8'b11000110;	//**   **
			16'h0573: data = 8'b11000110;	//**   **
			16'h0574: data = 8'b11000110;	//**   **
			16'h0575: data = 8'b11000110;	//**   **
			16'h0576: data = 8'b11000110;	//**   **
			16'h0577: data = 8'b11000110;	//**   **
			16'h0578: data = 8'b11010110;	//** * **
			16'h0579: data = 8'b11111110;	//*******
			16'h057a: data = 8'b11101110;	//*** ***  
			16'h057b: data = 8'b11000110;	//**   **
			16'h057c: data = 8'b00000000;	//
			16'h057d: data = 8'b00000000;	//
			16'h057e: data = 8'b00000000;	//
			16'h057f: data = 8'b00000000;	//
			// code x0058 (X)
			16'h0580: data = 8'b00000000;	//
			16'h0581: data = 8'b00000000;	//
			16'h0582: data = 8'b11000110;	//**   **
			16'h0583: data = 8'b11000110;	//**   **
			16'h0584: data = 8'b01101100;	// ** ** 
			16'h0585: data = 8'b00111000;	//  ***
			16'h0586: data = 8'b00111000;	//  *** 
			16'h0587: data = 8'b00111000;	//  ***
			16'h0588: data = 8'b00111000;	//  ***
			16'h0589: data = 8'b01101100;	// ** **
			16'h058a: data = 8'b11000110;	//**   **  
			16'h058b: data = 8'b11000110;	//**   **
			16'h058c: data = 8'b00000000;	//
			16'h058d: data = 8'b00000000;	//
			16'h058e: data = 8'b00000000;	//
			16'h058f: data = 8'b00000000;	//
			// code x0059 (Y)
			16'h0590: data = 8'b00000000;	//
			16'h0591: data = 8'b00000000;	//
			16'h0592: data = 8'b11000110;	//**   **
			16'h0593: data = 8'b11000110;	//**   **
			16'h0594: data = 8'b01101100;	// ** ** 
			16'h0595: data = 8'b00111000;	//  ***
			16'h0596: data = 8'b00011000;	//   ** 
			16'h0597: data = 8'b00011000;	//   **
			16'h0598: data = 8'b00011000;	//   **
			16'h0599: data = 8'b00011000;	//   **
			16'h059a: data = 8'b00011000;	//   **  
			16'h059b: data = 8'b00011000;	//   **
			16'h059c: data = 8'b00000000;	//
			16'h059d: data = 8'b00000000;	//
			16'h059e: data = 8'b00000000;	//
			16'h059f: data = 8'b00000000;	//
			// code x005a (Z)
			16'h05a0: data = 8'b00000000;	//
			16'h05a1: data = 8'b00000000;	//
			16'h05a2: data = 8'b11111110;	//*******
			16'h05a3: data = 8'b11111110;	//*******
			16'h05a4: data = 8'b00000110;	//     **  
			16'h05a5: data = 8'b00001100;	//    **
			16'h05a6: data = 8'b00011000;	//   ** 
			16'h05a7: data = 8'b00110000;	//  **
			16'h05a8: data = 8'b01100000;	// **
			16'h05a9: data = 8'b11000000;	//**
			16'h05aa: data = 8'b11111110;	//*******  
			16'h05ab: data = 8'b11111110;	//*******
			16'h05ac: data = 8'b00000000;	//
			16'h05ad: data = 8'b00000000;	//
			16'h05ae: data = 8'b00000000;	//
			16'h05af: data = 8'b00000000;	//
			// code x005b ([)
			16'h05b0: data = 8'b00000000;	//
			16'h05b1: data = 8'b00000000;	//
			16'h05b2: data = 8'b00000000;	//
			16'h05b3: data = 8'b00000000;	//
			16'h05b4: data = 8'b00000000;	//
			16'h05b5: data = 8'b00000000;	//
			16'h05b6: data = 8'b00000000;	//
			16'h05b7: data = 8'b00000000;	//
			16'h05b8: data = 8'b00000000;	//
			16'h05b9: data = 8'b00000000;	//
			16'h05ba: data = 8'b00000000;	//
			16'h05bb: data = 8'b00000000;	//
			16'h05bc: data = 8'b00000000;	//
			16'h05bd: data = 8'b00000000;	//
			16'h05be: data = 8'b00000000;	//
			16'h05bf: data = 8'b00000000;	//
			// code x005c (\)
			16'h05c0: data = 8'b00000000;	//
			16'h05c1: data = 8'b00000000;	//
			16'h05c2: data = 8'b00000000;	//
			16'h05c3: data = 8'b00000000;	//
			16'h05c4: data = 8'b00000000;	//
			16'h05c5: data = 8'b00000000;	//
			16'h05c6: data = 8'b00000000;	//
			16'h05c7: data = 8'b00000000;	//
			16'h05c8: data = 8'b00000000;	//
			16'h05c9: data = 8'b00000000;	//
			16'h05ca: data = 8'b00000000;	//
			16'h05cb: data = 8'b00000000;	//
			16'h05cc: data = 8'b00000000;	//
			16'h05cd: data = 8'b00000000;	//
			16'h05ce: data = 8'b00000000;	//
			16'h05cf: data = 8'b00000000;	//
			// code x005d (])
			16'h05d0: data = 8'b00000000;	//
			16'h05d1: data = 8'b00000000;	//
			16'h05d2: data = 8'b00000000;	//
			16'h05d3: data = 8'b00000000;	//
			16'h05d4: data = 8'b00000000;	//
			16'h05d5: data = 8'b00000000;	//
			16'h05d6: data = 8'b00000000;	//
			16'h05d7: data = 8'b00000000;	//
			16'h05d8: data = 8'b00000000;	//
			16'h05d9: data = 8'b00000000;	//
			16'h05da: data = 8'b00000000;	//
			16'h05db: data = 8'b00000000;	//
			16'h05dc: data = 8'b00000000;	//
			16'h05dd: data = 8'b00000000;	//
			16'h05de: data = 8'b00000000;	//
			16'h05df: data = 8'b00000000;	//
			// code x005e (^)
			16'h05e0: data = 8'b00000000;	//
			16'h05e1: data = 8'b00000000;	//
			16'h05e2: data = 8'b00000000;	//
			16'h05e3: data = 8'b00000000;	//
			16'h05e4: data = 8'b00000000;	//
			16'h05e5: data = 8'b00000000;	//
			16'h05e6: data = 8'b00000000;	//
			16'h05e7: data = 8'b00000000;	//
			16'h05e8: data = 8'b00000000;	//
			16'h05e9: data = 8'b00000000;	//
			16'h05ea: data = 8'b00000000;	//
			16'h05eb: data = 8'b00000000;	//
			16'h05ec: data = 8'b00000000;	//
			16'h05ed: data = 8'b00000000;	//
			16'h05ee: data = 8'b00000000;	//
			16'h05ef: data = 8'b00000000;	//
			// code x005f (_)
			16'h05f0: data = 8'b00000000;	//
			16'h05f1: data = 8'b00000000;	//
			16'h05f2: data = 8'b00000000;	//
			16'h05f3: data = 8'b00000000;	//
			16'h05f4: data = 8'b00000000;	//
			16'h05f5: data = 8'b00000000;	//
			16'h05f6: data = 8'b00000000;	//
			16'h05f7: data = 8'b00000000;	//
			16'h05f8: data = 8'b00000000;	//
			16'h05f9: data = 8'b00000000;	//
			16'h05fa: data = 8'b00000000;	//
			16'h05fb: data = 8'b00000000;	//
			16'h05fc: data = 8'b00000000;	//
			16'h05fd: data = 8'b00000000;	//
			16'h05fe: data = 8'b00000000;	//
			16'h05ff: data = 8'b00000000;	//
			// code x0060 (`)
			16'h0600: data = 8'b00000000;	//
			16'h0601: data = 8'b00000000;	//
			16'h0602: data = 8'b00000000;	//
			16'h0603: data = 8'b00000000;	//
			16'h0604: data = 8'b00000000;	//
			16'h0605: data = 8'b00000000;	//
			16'h0606: data = 8'b00000000;	//
			16'h0607: data = 8'b00000000;	//
			16'h0608: data = 8'b00000000;	//
			16'h0609: data = 8'b00000000;	//
			16'h060a: data = 8'b00000000;	//
			16'h060b: data = 8'b00000000;	//
			16'h060c: data = 8'b00000000;	//
			16'h060d: data = 8'b00000000;	//
			16'h060e: data = 8'b00000000;	//
			16'h060f: data = 8'b00000000;	//
			// code x0061 (a)
			16'h0610: data = 8'b00000000;	//
			16'h0611: data = 8'b00000000;	//
			16'h0612: data = 8'b00000000;	//
			16'h0613: data = 8'b00000000;	//
			16'h0614: data = 8'b00000000;	//
			16'h0615: data = 8'b00110110;	//
			16'h0616: data = 8'b11001110;	//
			16'h0617: data = 8'b11000110;	//
			16'h0618: data = 8'b11000110;	//
			16'h0619: data = 8'b11000110;	//
			16'h061a: data = 8'b01101110;	//
			16'h061b: data = 8'b00110110;	//
			16'h061c: data = 8'b00000000;	//
			16'h061d: data = 8'b00000000;	//
			16'h061e: data = 8'b00000000;	//
			16'h061f: data = 8'b00000000;	//
			// code x0062 (b)
			16'h0620: data = 8'b00000000;	//
			16'h0621: data = 8'b00000000;	//
			16'h0622: data = 8'b11000000;	//
			16'h0623: data = 8'b11000000;	//
			16'h0624: data = 8'b11000000;	//
			16'h0625: data = 8'b11011000;	//
			16'h0626: data = 8'b11101100;	//
			16'h0627: data = 8'b11000110;	//
			16'h0628: data = 8'b11000110;	//
			16'h0629: data = 8'b11000110;	//
			16'h062a: data = 8'b11101100;	//
			16'h062b: data = 8'b11011000;	//
			16'h062c: data = 8'b00000000;	//
			16'h062d: data = 8'b00000000;	//
			16'h062e: data = 8'b00000000;	//
			16'h062f: data = 8'b00000000;	//
			// code x0063 (c)
			16'h0630: data = 8'b00000000;	//
			16'h0631: data = 8'b00000000;	//
			16'h0632: data = 8'b00000000;	//
			16'h0633: data = 8'b00000000;	//
			16'h0634: data = 8'b00000000;	//
			16'h0635: data = 8'b00111000;	//
			16'h0636: data = 8'b01101100;	//
			16'h0637: data = 8'b11000110;	//
			16'h0638: data = 8'b11000000;	//
			16'h0639: data = 8'b11000110;	//
			16'h063a: data = 8'b01101100;	//
			16'h063b: data = 8'b00111000;	//
			16'h063c: data = 8'b00000000;	//
			16'h063d: data = 8'b00000000;	//
			16'h063e: data = 8'b00000000;	//
			16'h063f: data = 8'b00000000;	//
			// code x0064 (d)
			16'h0640: data = 8'b00000000;	//
			16'h0641: data = 8'b00000000;	//
			16'h0642: data = 8'b00000110;	//
			16'h0643: data = 8'b00000110;	//
			16'h0644: data = 8'b00000110;	//
			16'h0645: data = 8'b00110110;	//
			16'h0646: data = 8'b01101110;	//
			16'h0647: data = 8'b11000110;	//
			16'h0648: data = 8'b11000110;	//
			16'h0649: data = 8'b11000110;	//
			16'h064a: data = 8'b01101110;	//
			16'h064b: data = 8'b00110110;	//
			16'h064c: data = 8'b00000000;	//
			16'h064d: data = 8'b00000000;	//
			16'h064e: data = 8'b00000000;	//
			16'h064f: data = 8'b00000000;	//
			// code x0065 (e)
			16'h0650: data = 8'b00000000;	//
			16'h0651: data = 8'b00000000;	//
			16'h0652: data = 8'b00000000;	//
			16'h0653: data = 8'b00000000;	//
			16'h0654: data = 8'b00000000;	//
			16'h0655: data = 8'b00111000;	//
			16'h0656: data = 8'b01101100;	//
			16'h0657: data = 8'b11000110;	//
			16'h0658: data = 8'b11111110;	//
			16'h0659: data = 8'b11000000;	//
			16'h065a: data = 8'b01100110;	//
			16'h065b: data = 8'b00111100;	//
			16'h065c: data = 8'b00000000;	//
			16'h065d: data = 8'b00000000;	//
			16'h065e: data = 8'b00000000;	//
			16'h065f: data = 8'b00000000;	//
			// code x0066 (f)
			16'h0660: data = 8'b00000000;	//
			16'h0661: data = 8'b00000000;	//
			16'h0662: data = 8'b00111000;	//
			16'h0663: data = 8'b01101100;	//
			16'h0664: data = 8'b01100110;	//
			16'h0665: data = 8'b01100000;	//
			16'h0666: data = 8'b01100000;	//
			16'h0667: data = 8'b11111110;	//
			16'h0668: data = 8'b01100000;	//
			16'h0669: data = 8'b01100000;	//
			16'h066a: data = 8'b01100000;	//
			16'h066b: data = 8'b01100000;	//
			16'h066c: data = 8'b00000000;	//
			16'h066d: data = 8'b00000000;	//
			16'h066e: data = 8'b00000000;	//
			16'h066f: data = 8'b00000000;	//
			// code x0067 (g)
			16'h0670: data = 8'b00000000;	//
			16'h0671: data = 8'b00000000;	//
			16'h0672: data = 8'b00000000;	//
			16'h0673: data = 8'b00000000;	//
			16'h0674: data = 8'b00000000;	//
			16'h0675: data = 8'b00111011;	//-
			16'h0676: data = 8'b01000110;	//
			16'h0677: data = 8'b11000110;	//
			16'h0678: data = 8'b11000110;	//
			16'h0679: data = 8'b11000110;	//
			16'h067a: data = 8'b01000110;	//
			16'h067b: data = 8'b00111100;	//-
			16'h067c: data = 8'b00000110;	//
			16'h067d: data = 8'b11000110;	//
			16'h067e: data = 8'b00111000;	//-
			16'h067f: data = 8'b00000000;	//
			// code x0068 (h)
			16'h0680: data = 8'b00000000;	//
			16'h0681: data = 8'b00000000;	//
			16'h0682: data = 8'b11000000;	//-
			16'h0683: data = 8'b11000000;	//
			16'h0684: data = 8'b11000000;	//
			16'h0685: data = 8'b11111100;	//-
			16'h0686: data = 8'b11000110;	//
			16'h0687: data = 8'b11000110;	//
			16'h0688: data = 8'b11000110;	//
			16'h0689: data = 8'b11000110;	//
			16'h068a: data = 8'b11000110;	//
			16'h068b: data = 8'b11000110;	//-
			16'h068c: data = 8'b00000000;	//
			16'h068d: data = 8'b00000000;	//
			16'h068e: data = 8'b00000000;	//
			16'h068f: data = 8'b00000000;	//
			// code x0069 (i)
			16'h0690: data = 8'b00000000;	//
			16'h0691: data = 8'b00000000;	//
			16'h0692: data = 8'b00011000;	//
			16'h0693: data = 8'b00011000;	//
			16'h0694: data = 8'b00000000;	//
			16'h0695: data = 8'b01111000;	//-
			16'h0696: data = 8'b00011000;	//
			16'h0697: data = 8'b00011000;	//
			16'h0698: data = 8'b00011000;	//
			16'h0699: data = 8'b00011000;	//
			16'h069a: data = 8'b00011000;	//
			16'h069b: data = 8'b11111110;	//
			16'h069c: data = 8'b00000000;	//
			16'h069d: data = 8'b00000000;	//-
			16'h069e: data = 8'b00000000;	//
			16'h069f: data = 8'b00000000;	//
			// code x006a (j)
			16'h06a0: data = 8'b00000000;	//
			16'h06a1: data = 8'b00000000;	//
			16'h06a2: data = 8'b00011000;	//
			16'h06a3: data = 8'b00011000;	//
			16'h06a4: data = 8'b00000000;	//
			16'h06a5: data = 8'b00111100;	//-
			16'h06a6: data = 8'b00001100;	//
			16'h06a7: data = 8'b00001100;	//
			16'h06a8: data = 8'b00001100;	//
			16'h06a9: data = 8'b00001100;	//
			16'h06aa: data = 8'b00001100;	//
			16'h06ab: data = 8'b00001100;	//-
			16'h06ac: data = 8'b00001100;	//
			16'h06ad: data = 8'b11001100;	//
			16'h06ae: data = 8'b01111000;	//
			16'h06af: data = 8'b00000000;	//
			// code x006b (k)
			16'h06b0: data = 8'b00000000;	//
			16'h06b1: data = 8'b00000000;	//
			16'h06b2: data = 8'b11000000;	//-
			16'h06b3: data = 8'b11000000;	//-
			16'h06b4: data = 8'b11000000;	//-
			16'h06b5: data = 8'b11000110;	//x
			16'h06b6: data = 8'b11001100;	//x
			16'h06b7: data = 8'b11010000;	//x
			16'h06b8: data = 8'b11100000;	//x
			16'h06b9: data = 8'b11010000;	//x
			16'h06ba: data = 8'b11001100;	//x
			16'h06bb: data = 8'b11000110;	//x
			16'h06bc: data = 8'b00000000;	//-
			16'h06bd: data = 8'b00000000;	//-
			16'h06be: data = 8'b00000000;	//-
			16'h06bf: data = 8'b00000000;	//
			// code x006c (l)
			16'h06c0: data = 8'b00000000;	//
			16'h06c1: data = 8'b00000000;	//
			16'h06c2: data = 8'b01100000;	//-
			16'h06c3: data = 8'b01100000;	//-
			16'h06c4: data = 8'b01100000;	//-
			16'h06c5: data = 8'b01100000;	//x
			16'h06c6: data = 8'b01100000;	//x
			16'h06c7: data = 8'b01100000;	//x
			16'h06c8: data = 8'b01100000;	//x
			16'h06c9: data = 8'b01100000;	//x
			16'h06ca: data = 8'b01100000;	//x
			16'h06cb: data = 8'b00111100;	//x
			16'h06cc: data = 8'b00000000;	//-
			16'h06cd: data = 8'b00000000;	//-
			16'h06ce: data = 8'b00000000;	//-
			16'h06cf: data = 8'b00000000;	//
			// code x006d (m)
			16'h06d0: data = 8'b00000000;	//
			16'h06d1: data = 8'b00000000;	//
			16'h06d2: data = 8'b00000000;	//-
			16'h06d3: data = 8'b00000000;	//-
			16'h06d4: data = 8'b00000000;	//-
			16'h06d5: data = 8'b11101100;	//x
			16'h06d6: data = 8'b11010110;	//x
			16'h06d7: data = 8'b11010110;	//x
			16'h06d8: data = 8'b11010110;	//x
			16'h06d9: data = 8'b11010110;	//x
			16'h06da: data = 8'b11010110;	//x
			16'h06db: data = 8'b11000110;	//x
			16'h06dc: data = 8'b00000000;	//-
			16'h06dd: data = 8'b00000000;	//-
			16'h06de: data = 8'b00000000;	//-
			16'h06df: data = 8'b00000000;	//
			// code x006e (n)
			16'h06e0: data = 8'b00000000;	//
			16'h06e1: data = 8'b00000000;	//
			16'h06e2: data = 8'b00000000;	//-
			16'h06e3: data = 8'b00000000;	//-
			16'h06e4: data = 8'b00000000;	//-
			16'h06e5: data = 8'b10111100;	//x
			16'h06e6: data = 8'b11000110;	//x
			16'h06e7: data = 8'b11000110;	//x
			16'h06e8: data = 8'b11000110;	//x
			16'h06e9: data = 8'b11000110;	//x
			16'h06ea: data = 8'b11000110;	//x
			16'h06eb: data = 8'b11000110;	//x
			16'h06ec: data = 8'b00000000;	//-
			16'h06ed: data = 8'b00000000;	//-
			16'h06ee: data = 8'b00000000;	//-
			16'h06ef: data = 8'b00000000;	//
			// code x006f (o)
			16'h06f0: data = 8'b00000000;	//
			16'h06f1: data = 8'b00000000;	//
			16'h06f2: data = 8'b00000000;	//-
			16'h06f3: data = 8'b00000000;	//-
			16'h06f4: data = 8'b00000000;	//-
			16'h06f5: data = 8'b01111100;	//x
			16'h06f6: data = 8'b11000110;	//x
			16'h06f7: data = 8'b11000110;	//x
			16'h06f8: data = 8'b11000110;	//x
			16'h06f9: data = 8'b11000110;	//x
			16'h06fa: data = 8'b11000110;	//x
			16'h06fb: data = 8'b01111100;	//x
			16'h06fc: data = 8'b00000000;	//-
			16'h06fd: data = 8'b00000000;	//-
			16'h06fe: data = 8'b00000000;	//-
			16'h06ff: data = 8'b00000000;	//
			// code x0070 (p)
			16'h0700: data = 8'b00000000;	//
			16'h0701: data = 8'b00000000;	//
			16'h0702: data = 8'b00000000;	//-
			16'h0703: data = 8'b00000000;	//-
			16'h0704: data = 8'b00000000;	//-
			16'h0705: data = 8'b11111100;	//x
			16'h0706: data = 8'b11000110;	//x
			16'h0707: data = 8'b11000110;	//x
			16'h0708: data = 8'b11000110;	//x
			16'h0709: data = 8'b11000110;	//x
			16'h070a: data = 8'b11000110;	//x
			16'h070b: data = 8'b11111100;	//x
			16'h070c: data = 8'b11000000;	//-
			16'h070d: data = 8'b11000000;	//-
			16'h070e: data = 8'b11000000;	//-
			16'h070f: data = 8'b00000000;	//
			// code x0071 (q)
			16'h0710: data = 8'b00000000;	//
			16'h0711: data = 8'b00000000;	//
			16'h0712: data = 8'b00000000;	//-
			16'h0713: data = 8'b00000000;	//-
			16'h0714: data = 8'b00000000;	//-
			16'h0715: data = 8'b01111110;	//x
			16'h0716: data = 8'b11000110;	//x
			16'h0717: data = 8'b11000110;	//x
			16'h0718: data = 8'b11000110;	//x
			16'h0719: data = 8'b11000110;	//x
			16'h071a: data = 8'b11000110;	//x
			16'h071b: data = 8'b01111110;	//x
			16'h071c: data = 8'b00000110;	//-
			16'h071d: data = 8'b00000110;	//-
			16'h071e: data = 8'b00000110;	//-
			16'h071f: data = 8'b00000000;	//
			// code x0072 (r)
			16'h0720: data = 8'b00000000;	//
			16'h0721: data = 8'b00000000;	//
			16'h0722: data = 8'b00000000;	//-
			16'h0723: data = 8'b00000000;	//-
			16'h0724: data = 8'b00000000;	//-
			16'h0725: data = 8'b10111100;	//x
			16'h0726: data = 8'b11000010;	//x
			16'h0727: data = 8'b11000000;	//x
			16'h0728: data = 8'b11000000;	//x
			16'h0729: data = 8'b11000000;	//x
			16'h072a: data = 8'b11000000;	//x
			16'h072b: data = 8'b11000000;	//x
			16'h072c: data = 8'b00000000;	//-
			16'h072d: data = 8'b00000000;	//-
			16'h072e: data = 8'b00000000;	//-
			16'h072f: data = 8'b00000000;	//
			// code x0073 (s)
			16'h0730: data = 8'b00000000;	//
			16'h0731: data = 8'b00000000;	//
			16'h0732: data = 8'b00000000;	//-
			16'h0733: data = 8'b00000000;	//-
			16'h0734: data = 8'b00000000;	//-
			16'h0735: data = 8'b01111110;	//x
			16'h0736: data = 8'b11000000;	//x
			16'h0737: data = 8'b11000000;	//x
			16'h0738: data = 8'b01111100;	//x
			16'h0739: data = 8'b00000110;	//x
			16'h073a: data = 8'b00000110;	//x
			16'h073b: data = 8'b11111100;	//x
			16'h073c: data = 8'b00000000;	//-
			16'h073d: data = 8'b00000000;	//-
			16'h073e: data = 8'b00000000;	//-
			16'h073f: data = 8'b00000000;	//
			// code x0074 (t)
			16'h0740: data = 8'b00000000;	//
			16'h0741: data = 8'b00000000;	//
			16'h0742: data = 8'b11000000;	//-
			16'h0743: data = 8'b11000000;	//-
			16'h0744: data = 8'b11000000;	//-
			16'h0745: data = 8'b11000000;	//x
			16'h0746: data = 8'b11111000;	//x
			16'h0747: data = 8'b11100000;	//x
			16'h0748: data = 8'b11000000;	//x
			16'h0749: data = 8'b11000110;	//x
			16'h074a: data = 8'b11000110;	//x
			16'h074b: data = 8'b01111100;	//x
			16'h074c: data = 8'b00000000;	//-
			16'h074d: data = 8'b00000000;	//-
			16'h074e: data = 8'b00000000;	//-
			16'h074f: data = 8'b00000000;	//
			// code x0075 (u)
			16'h0750: data = 8'b00000000;	//
			16'h0751: data = 8'b00000000;	//
			16'h0752: data = 8'b00000000;	//-
			16'h0753: data = 8'b00000000;	//-
			16'h0754: data = 8'b00000000;	//-
			16'h0755: data = 8'b11000110;	//x
			16'h0756: data = 8'b11000110;	//x
			16'h0757: data = 8'b11000110;	//x
			16'h0758: data = 8'b11000110;	//x
			16'h0759: data = 8'b11000110;	//x
			16'h075a: data = 8'b11000110;	//x
			16'h075b: data = 8'b00111010;	//x
			16'h075c: data = 8'b00000000;	//-
			16'h075d: data = 8'b00000000;	//-
			16'h075e: data = 8'b00000000;	//-
			16'h075f: data = 8'b00000000;	//
			// code x0076 (v)
			16'h0760: data = 8'b00000000;	//
			16'h0761: data = 8'b00000000;	//
			16'h0762: data = 8'b00000000;	//-
			16'h0763: data = 8'b00000000;	//-
			16'h0764: data = 8'b00000000;	//-
			16'h0765: data = 8'b11000110;	//x
			16'h0766: data = 8'b11000110;	//x
			16'h0767: data = 8'b11000110;	//x
			16'h0768: data = 8'b11000110;	//x
			16'h0769: data = 8'b01000100;	//x
			16'h076a: data = 8'b00101000;	//x
			16'h076b: data = 8'b00010000;	//x
			16'h076c: data = 8'b00000000;	//-
			16'h076d: data = 8'b00000000;	//-
			16'h076e: data = 8'b00000000;	//-
			16'h076f: data = 8'b00000000;	//
			// code x0077 (w)
			16'h0770: data = 8'b00000000;	//
			16'h0771: data = 8'b00000000;	//
			16'h0772: data = 8'b00000000;	//-
			16'h0773: data = 8'b00000000;	//-
			16'h0774: data = 8'b00000000;	//-
			16'h0775: data = 8'b11000010;	//x
			16'h0776: data = 8'b11000010;	//x
			16'h0777: data = 8'b11011010;	//x
			16'h0778: data = 8'b11011010;	//x
			16'h0779: data = 8'b11011010;	//x
			16'h077a: data = 8'b01100110;	//x
			16'h077b: data = 8'b01000100;	//x
			16'h077c: data = 8'b00000000;	//-
			16'h077d: data = 8'b00000000;	//-
			16'h077e: data = 8'b00000000;	//-
			16'h077f: data = 8'b00000000;	//
			// code x0078 (x)
			16'h0780: data = 8'b00000000;	//
			16'h0781: data = 8'b00000000;	//
			16'h0782: data = 8'b00000000;	//-
			16'h0783: data = 8'b00000000;	//-
			16'h0784: data = 8'b00000000;	//-
			16'h0785: data = 8'b11000110;	//x
			16'h0786: data = 8'b11000110;	//x
			16'h0787: data = 8'b01101100;	//x
			16'h0788: data = 8'b00010000;	//x
			16'h0789: data = 8'b01101100;	//x
			16'h078a: data = 8'b11000110;	//x
			16'h078b: data = 8'b11000110;	//x
			16'h078c: data = 8'b00000000;	//-
			16'h078d: data = 8'b00000000;	//-
			16'h078e: data = 8'b00000000;	//-
			16'h078f: data = 8'b00000000;	//
			// code x0079 (y)
			16'h0790: data = 8'b00000000;	//
			16'h0791: data = 8'b00000000;	//
			16'h0792: data = 8'b00000000;	//-
			16'h0793: data = 8'b00000000;	//-
			16'h0794: data = 8'b00000000;	//-
			16'h0795: data = 8'b11000110;	//x
			16'h0796: data = 8'b11000110;	//x
			16'h0797: data = 8'b11000110;	//x
			16'h0798: data = 8'b11000110;	//x
			16'h0799: data = 8'b11000110;	//x
			16'h079a: data = 8'b01000110;	//x
			16'h079b: data = 8'b00111110;	//x
			16'h079c: data = 8'b00000110;	//-
			16'h079d: data = 8'b01000110;	//-
			16'h079e: data = 8'b00111110;	//-
			16'h079f: data = 8'b00000000;	//
			// code x007a (z)
			16'h07a0: data = 8'b00000000;	//
			16'h07a1: data = 8'b00000000;	//
			16'h07a2: data = 8'b00000000;	//-
			16'h07a3: data = 8'b00000000;	//-
			16'h07a4: data = 8'b00000000;	//-
			16'h07a5: data = 8'b11111110;	//x
			16'h07a6: data = 8'b00000110;	//x
			16'h07a7: data = 8'b00001100;	//x
			16'h07a8: data = 8'b00011000;	//x
			16'h07a9: data = 8'b00110000;	//x
			16'h07aa: data = 8'b01100000;	//x
			16'h07ab: data = 8'b11111110;	//x
			16'h07ac: data = 8'b00000000;	//-
			16'h07ad: data = 8'b00000000;	//-
			16'h07ae: data = 8'b00000000;	//-
			16'h07af: data = 8'b00000000;	//
			// code x007b ({)
			16'h07b0: data = 8'b00000000;	//
			16'h07b1: data = 8'b00000000;	//
			16'h07b2: data = 8'b00000000;	//
			16'h07b3: data = 8'b00000000;	//
			16'h07b4: data = 8'b00000000;	//
			16'h07b5: data = 8'b00000000;	//
			16'h07b6: data = 8'b00000000;	//
			16'h07b7: data = 8'b00000000;	//
			16'h07b8: data = 8'b00000000;	//
			16'h07b9: data = 8'b00000000;	//
			16'h07ba: data = 8'b00000000;	//
			16'h07bb: data = 8'b00000000;	//
			16'h07bc: data = 8'b00000000;	//
			16'h07bd: data = 8'b00000000;	//
			16'h07be: data = 8'b00000000;	//
			16'h07bf: data = 8'b00000000;	//
			// code x007c (|)
			16'h07c0: data = 8'b00000000;	//
			16'h07c1: data = 8'b00000000;	//
			16'h07c2: data = 8'b00010000;	//   *
			16'h07c3: data = 8'b00010000;	//   *
			16'h07c4: data = 8'b00010000;	//   *
			16'h07c5: data = 8'b00010000;	//   *
			16'h07c6: data = 8'b00010000;	//   *
			16'h07c7: data = 8'b00010000;	//   *
			16'h07c8: data = 8'b00010000;	//   *
			16'h07c9: data = 8'b00010000;	//   *
			16'h07ca: data = 8'b00010000;	//   *
			16'h07cb: data = 8'b00010000;	//   *
			16'h07cc: data = 8'b00000000;	//
			16'h07cd: data = 8'b00000000;	//
			16'h07ce: data = 8'b00000000;	//
			16'h07cf: data = 8'b00000000;	//
			// code x007d (})
			16'h07d0: data = 8'b00000000;	//
			16'h07d1: data = 8'b00000000;	//
			16'h07d2: data = 8'b00000000;	//
			16'h07d3: data = 8'b00000000;	//
			16'h07d4: data = 8'b00000000;	//
			16'h07d5: data = 8'b00000000;	//
			16'h07d6: data = 8'b00000000;	//
			16'h07d7: data = 8'b00000000;	//
			16'h07d8: data = 8'b00000000;	//
			16'h07d9: data = 8'b00000000;	//
			16'h07da: data = 8'b00000000;	//
			16'h07db: data = 8'b00000000;	//
			16'h07dc: data = 8'b00000000;	//
			16'h07dd: data = 8'b00000000;	//
			16'h07de: data = 8'b00000000;	//
			16'h07df: data = 8'b00000000;	//
			// code x007e (~)
			16'h07e0: data = 8'b00000000;	//
			16'h07e1: data = 8'b00000000;	//
			16'h07e2: data = 8'b00000000;	//
			16'h07e3: data = 8'b00000000;	//
			16'h07e4: data = 8'b00000000;	//
			16'h07e5: data = 8'b00000000;	//
			16'h07e6: data = 8'b00000000;	//
			16'h07e7: data = 8'b00000000;	//
			16'h07e8: data = 8'b00000000;	//
			16'h07e9: data = 8'b00000000;	//
			16'h07ea: data = 8'b00000000;	//
			16'h07eb: data = 8'b00000000;	//
			16'h07ec: data = 8'b00000000;	//
			16'h07ed: data = 8'b00000000;	//
			16'h07ee: data = 8'b00000000;	//
			16'h07ef: data = 8'b00000000;	//
			// code x007f (del) delete, which is the all-one pattern
			16'h07f0: data = 8'b11111111;	//********
			16'h07f1: data = 8'b11111111;	//********
			16'h07f2: data = 8'b11111111;	//********
			16'h07f3: data = 8'b11111111;	//********
			16'h07f4: data = 8'b11111111;	//********
			16'h07f5: data = 8'b11111111;	//********
			16'h07f6: data = 8'b11111111;	//********
			16'h07f7: data = 8'b11111111;	//********
			16'h07f8: data = 8'b11111111;	//********
			16'h07f9: data = 8'b11111111;	//********
			16'h07fa: data = 8'b11111111;	//********
			16'h07fb: data = 8'b11111111;	//********
			16'h07fc: data = 8'b11111111;	//********
			16'h07fd: data = 8'b11111111;	//********
			16'h07fe: data = 8'b11111111;	//********
			16'h07ff: data = 8'b11111111;	//********
			
			// code xB881 (korkai)
            16'h8810: data = 8'b00000000;	//
            16'h8811: data = 8'b00000000;	//
            16'h8812: data = 8'b00000000;	//
            16'h8813: data = 8'b00000000;	//
            16'h8814: data = 8'b00000000;	//
            16'h8815: data = 8'b00111000;	//
            16'h8816: data = 8'b01101100;	//
            16'h8817: data = 8'b11000110;	//
            16'h8818: data = 8'b01100110;	//
            16'h8819: data = 8'b11000110;	//
            16'h881a: data = 8'b11000110;	//
            16'h881b: data = 8'b11000110;	//
            16'h881c: data = 8'b00000000;	//
            16'h881d: data = 8'b00000000;	//
            16'h881e: data = 8'b00000000;	//
            16'h881f: data = 8'b00000000;	//
            
            // code xB882 (khor-kai)
            16'h8820: data = 8'b00000000;
            16'h8821: data = 8'b00000000;
            16'h8822: data = 8'b00000000;
            16'h8823: data = 8'b00000000;
            16'h8824: data = 8'b00000000;
            16'h8825: data = 8'b11000110;
            16'h8826: data = 8'b10100110;
            16'h8827: data = 8'b01100110;
            16'h8828: data = 8'b11000110;
            16'h8829: data = 8'b11000110;
            16'h882A: data = 8'b01101100;
            16'h882B: data = 8'b00111000;
            16'h882C: data = 8'b00000000;
            16'h882D: data = 8'b00000000;
            16'h882E: data = 8'b00000000;
            16'h882F: data = 8'b00000000;
            
            // code xB883 (khor-kood)
            16'h8830: data = 8'b00000000;
            16'h8831: data = 8'b00000000;
            16'h8832: data = 8'b00000000;
            16'h8833: data = 8'b00000000;
            16'h8834: data = 8'b00000000;
            16'h8835: data = 8'b01010110;
            16'h8836: data = 8'b10110110;
            16'h8837: data = 8'b01100110;
            16'h8838: data = 8'b11000110;
            16'h8839: data = 8'b11000110;
            16'h883A: data = 8'b01101100;
            16'h883B: data = 8'b00111000;
            16'h883C: data = 8'b00000000;
            16'h883D: data = 8'b00000000;
            16'h883E: data = 8'b00000000;
            16'h883F: data = 8'b00000000;
            
            // code xB884 (buffalo)
            16'h8840: data = 8'b00000000;
            16'h8841: data = 8'b00000000;
            16'h8842: data = 8'b00000000;
            16'h8843: data = 8'b00000000;
            16'h8844: data = 8'b00000000;
            16'h8845: data = 8'b00111000;
            16'h8846: data = 8'b01101100;
            16'h8847: data = 8'b11000110;
            16'h8848: data = 8'b10110110;
            16'h8849: data = 8'b11101110;
            16'h884A: data = 8'b11111110;
            16'h884B: data = 8'b11000110;
            16'h884C: data = 8'b00000000;
            16'h884D: data = 8'b00000000;
            16'h884E: data = 8'b00000000;
            16'h884F: data = 8'b00000000;
            
            // code xB885 (human)
            16'h8850: data = 8'b00000000;
            16'h8851: data = 8'b00000000;
            16'h8852: data = 8'b00000000;
            16'h8853: data = 8'b00000000;
            16'h8854: data = 8'b00000000;
            16'h8855: data = 8'b00101000;
            16'h8856: data = 8'b01111100;
            16'h8857: data = 8'b11000110;
            16'h8858: data = 8'b10110110;
            16'h8859: data = 8'b11101110;
            16'h885A: data = 8'b11111110;
            16'h885B: data = 8'b11000110;
            16'h885C: data = 8'b00000000;
            16'h885D: data = 8'b00000000;
            16'h885E: data = 8'b00000000;
            16'h885F: data = 8'b00000000;
            
            // code xB886 (khor-bell)
            16'h8860: data = 8'b00000000;
            16'h8861: data = 8'b00000000;
            16'h8862: data = 8'b00000000;
            16'h8863: data = 8'b00000000;
            16'h8864: data = 8'b00000000;
            16'h8865: data = 8'b01010110;
            16'h8866: data = 8'b10110110;
            16'h8867: data = 8'b01100110;
            16'h8868: data = 8'b01100110;
            16'h8869: data = 8'b11100110;
            16'h886A: data = 8'b10111110;
            16'h886B: data = 8'b11101110;
            16'h886C: data = 8'b00000000;
            16'h886D: data = 8'b00000000;
            16'h886E: data = 8'b00000000;
            16'h886F: data = 8'b00000000;
            
            // code xB887 (ngor-ngu)
            16'h8870: data = 8'b00000000;	//
            16'h8871: data = 8'b00000000;	//
            16'h8872: data = 8'b00000000;	//
            16'h8873: data = 8'b00000000;	//
            16'h8874: data = 8'b00000000;	//
            16'h8875: data = 8'b00000110;	//
            16'h8876: data = 8'b00001010;	//
            16'h8877: data = 8'b00000110;	//
            16'h8878: data = 8'b11000110;	//
            16'h8879: data = 8'b01100110;	//
            16'h887a: data = 8'b00110110;	//
            16'h887b: data = 8'b00011100;	//
            16'h887c: data = 8'b00000000;	//
            16'h887d: data = 8'b00000000;	//
            16'h887e: data = 8'b00000000;	//
            16'h887f: data = 8'b00000000;	//
            
            // code xB888 (jor-jan)
            16'h8880: data = 8'b00000000;	//
            16'h8881: data = 8'b00000000;	//
            16'h8882: data = 8'b00000000;	//
            16'h8883: data = 8'b00000000;	//
            16'h8884: data = 8'b00000000;	//
            16'h8885: data = 8'b00111000;	//
            16'h8886: data = 8'b01101100;	//
            16'h8887: data = 8'b10000110;	//
            16'h8888: data = 8'b00100110;	//
            16'h8889: data = 8'b01010110;	//
            16'h888a: data = 8'b00110110;	//
            16'h888b: data = 8'b00001110;	//
            16'h888c: data = 8'b00000000;	//
            16'h888d: data = 8'b00000000;	//
            16'h888e: data = 8'b00000000;	//
            16'h888f: data = 8'b00000000;	//
            
            // code xB889 (chor-ching)
            16'h8890: data = 8'b00000000;
            16'h8891: data = 8'b00000000;
            16'h8892: data = 8'b00000000;
            16'h8893: data = 8'b00000000;
            16'h8894: data = 8'b00000000;
            16'h8895: data = 8'b01111000;
            16'h8896: data = 8'b10001100;
            16'h8897: data = 8'b01000110;
            16'h8898: data = 8'b10100110;
            16'h8899: data = 8'b11101110;
            16'h889A: data = 8'b01111010;
            16'h889B: data = 8'b01101100;
            16'h889C: data = 8'b00000000;
            16'h889D: data = 8'b00000000;
            16'h889E: data = 8'b00000000;
            16'h889F: data = 8'b00000000;
            
            // code xB88A (chor-chang)
            16'h88A0: data = 8'b00000000;
            16'h88A1: data = 8'b00000000;
            16'h88A2: data = 8'b00000000;
            16'h88A3: data = 8'b00000010;
            16'h88A4: data = 8'b00000010;
            16'h88A5: data = 8'b01000110;
            16'h88A6: data = 8'b10101100;
            16'h88A7: data = 8'b11100110;
            16'h88A8: data = 8'b01000110;
            16'h88A9: data = 8'b11000110;
            16'h88AA: data = 8'b01101100;
            16'h88AB: data = 8'b00111000;
            16'h88AC: data = 8'b00000000;
            16'h88AD: data = 8'b00000000;
            16'h88AE: data = 8'b00000000;
            16'h88AF: data = 8'b00000000;
            
            // code xB88B (zor-so)
            16'h88B0: data = 8'b00000000;
            16'h88B1: data = 8'b00000000;
            16'h88B2: data = 8'b00000000;
            16'h88B3: data = 8'b00000010;
            16'h88B4: data = 8'b00000010;
            16'h88B5: data = 8'b01010110;
            16'h88B6: data = 8'b10110100;
            16'h88B7: data = 8'b11100110;
            16'h88B8: data = 8'b01000110;
            16'h88B9: data = 8'b11100110;
            16'h88BA: data = 8'b01101100;
            16'h88BB: data = 8'b00111000;
            16'h88BC: data = 8'b00000000;
            16'h88BD: data = 8'b00000000;
            16'h88BE: data = 8'b00000000;
            16'h88BF: data = 8'b00000000;
            
            // code xB88C (chor-cher)
            16'h88C0: data = 8'b00000000;
            16'h88C1: data = 8'b00000000;
            16'h88C2: data = 8'b00000000;
            16'h88C3: data = 8'b00000000;
            16'h88C4: data = 8'b00000000;
            16'h88C5: data = 8'b01110010;
            16'h88C6: data = 8'b11010010;
            16'h88C7: data = 8'b01010010;
            16'h88C8: data = 8'b11011010;
            16'h88C9: data = 8'b11011110;
            16'h88CA: data = 8'b10101110;
            16'h88CB: data = 8'b01111110;
            16'h88CC: data = 8'b00000000;
            16'h88CD: data = 8'b00000000;
            16'h88CE: data = 8'b00000000;
            16'h88CF: data = 8'b00000000;
            
            // code xB88D (yor-ying)
            16'h88D0: data = 8'b00000000;
            16'h88D1: data = 8'b00000000;
            16'h88D2: data = 8'b00000000;
            16'h88D3: data = 8'b00000000;
            16'h88D4: data = 8'b00000000;
            16'h88D5: data = 8'b01111010;
            16'h88D6: data = 8'b11001010;
            16'h88D7: data = 8'b01001010;
            16'h88D8: data = 8'b11001010;
            16'h88D9: data = 8'b11101010;
            16'h88DA: data = 8'b10101110;
            16'h88DB: data = 8'b01101110;
            16'h88DC: data = 8'b00000000;
            16'h88DD: data = 8'b00001010;
            16'h88DE: data = 8'b00001110;
            16'h88DF: data = 8'b00000000;
            
            // code xB88E (tor-unknow-1)
            16'h88E0: data = 8'b00000000;
            16'h88E1: data = 8'b00000000;
            16'h88E2: data = 8'b00000000;
            16'h88E3: data = 8'b00000000;
            16'h88E4: data = 8'b00000000;
            16'h88E5: data = 8'b01111100;
            16'h88E6: data = 8'b11101110;
            16'h88E7: data = 8'b01000110;
            16'h88E8: data = 8'b01100110;
            16'h88E9: data = 8'b11100110;
            16'h88EA: data = 8'b10100110;
            16'h88EB: data = 8'b01100110;
            16'h88EC: data = 8'b00010110;
            16'h88ED: data = 8'b00101110;
            16'h88EE: data = 8'b00011110;
            16'h88EF: data = 8'b00000000;
            
            // code xB88F (tor-unknow-2)
            16'h88F0: data = 8'b00000000;
            16'h88F1: data = 8'b00000000;
            16'h88F2: data = 8'b00000000;
            16'h88F3: data = 8'b00000000;
            16'h88F4: data = 8'b00000000;
            16'h88F5: data = 8'b01111100;
            16'h88F6: data = 8'b11101110;
            16'h88F7: data = 8'b01000110;
            16'h88F8: data = 8'b01100110;
            16'h88F9: data = 8'b11100110;
            16'h88FA: data = 8'b10100110;
            16'h88FB: data = 8'b01100110;
            16'h88FC: data = 8'b00010110;
            16'h88FD: data = 8'b00101110;
            16'h88FE: data = 8'b00010110;
            16'h88FF: data = 8'b00000000;
            
            // code xB890 (thor-than)
            16'h8900: data = 8'b00000000;
            16'h8901: data = 8'b00000000;
            16'h8902: data = 8'b00000000;
            16'h8903: data = 8'b00000000;
            16'h8904: data = 8'b00000000;
            16'h8905: data = 8'b01111110;
            16'h8906: data = 8'b11100000;
            16'h8907: data = 8'b00111110;
            16'h8908: data = 8'b00010110;
            16'h8909: data = 8'b00101110;
            16'h890A: data = 8'b00011110;
            16'h890B: data = 8'b00000110;
            16'h890C: data = 8'b00100000;
            16'h890D: data = 8'b01010110;
            16'h890E: data = 8'b01101100;
            16'h890F: data = 8'b00000000;
            
            // code xB891 (thor-ngang-two)
            16'h8910: data = 8'b00000000;
            16'h8911: data = 8'b00000000;
            16'h8912: data = 8'b00000000;
            16'h8913: data = 8'b00000000;
            16'h8914: data = 8'b00000000;
            16'h8915: data = 8'b01010110;
            16'h8916: data = 8'b10100110;
            16'h8917: data = 8'b01101110;
            16'h8918: data = 8'b01111110;
            16'h8919: data = 8'b01110110;
            16'h891A: data = 8'b01100110;
            16'h891B: data = 8'b01100110;
            16'h891C: data = 8'b00000000;
            16'h891D: data = 8'b00000000;
            16'h891E: data = 8'b00000000;
            16'h891F: data = 8'b00000000;
            
            // code xB892 (thor-phu-thao)
            16'h8920: data = 8'b00000000;
            16'h8921: data = 8'b00000000;
            16'h8922: data = 8'b00000000;
            16'h8923: data = 8'b00000000;
            16'h8924: data = 8'b00000000;
            16'h8925: data = 8'b01010010;
            16'h8926: data = 8'b10101010;
            16'h8927: data = 8'b10001010;
            16'h8928: data = 8'b10110010;
            16'h8929: data = 8'b11101010;
            16'h892A: data = 8'b11011110;
            16'h892B: data = 8'b11010110;
            16'h892C: data = 8'b00000000;
            16'h892D: data = 8'b00000000;
            16'h892E: data = 8'b00000000;
            16'h892F: data = 8'b00000000;
            
            // code xB893 (nor-nen)
            16'h8930: data = 8'b00000000;
            16'h8931: data = 8'b00000000;
            16'h8932: data = 8'b00000000;
            16'h8933: data = 8'b00000000;
            16'h8934: data = 8'b00000000;
            16'h8935: data = 8'b01110010;
            16'h8936: data = 8'b11011010;
            16'h8937: data = 8'b10001010;
            16'h8938: data = 8'b10001010;
            16'h8939: data = 8'b11001110;
            16'h893A: data = 8'b10101010;
            16'h893B: data = 8'b01001010;
            16'h893C: data = 8'b00000000;
            16'h893D: data = 8'b00000000;
            16'h893E: data = 8'b00000000;
            16'h893F: data = 8'b00000000;
            
            // code xB894 (door-dek)
            16'h8940: data = 8'b00000000;
            16'h8941: data = 8'b00000000;
            16'h8942: data = 8'b00000000;
            16'h8943: data = 8'b00000000;
            16'h8944: data = 8'b00000000;
            16'h8945: data = 8'b00111000;
            16'h8946: data = 8'b01101100;
            16'h8947: data = 8'b11000110;
            16'h8948: data = 8'b10010010;
            16'h8949: data = 8'b10101010;
            16'h894A: data = 8'b11110010;
            16'h894B: data = 8'b11100010;
            16'h894C: data = 8'b00000000;
            16'h894D: data = 8'b00000000;
            16'h894E: data = 8'b00000000;
            16'h894F: data = 8'b00000000;
            
            // code xB895 (tor-tao)
            16'h8950: data = 8'b00000000;
            16'h8951: data = 8'b00000000;
            16'h8952: data = 8'b00000000;
            16'h8953: data = 8'b00000000;
            16'h8954: data = 8'b00000000;
            16'h8955: data = 8'b00101000;
            16'h8956: data = 8'b01111100;
            16'h8957: data = 8'b11000110;
            16'h8958: data = 8'b10010010;
            16'h8959: data = 8'b10101010;
            16'h895A: data = 8'b11110010;
            16'h895B: data = 8'b11100010;
            16'h895C: data = 8'b00000000;
            16'h895D: data = 8'b00000000;
            16'h895E: data = 8'b00000000;
            16'h895F: data = 8'b00000000;
            
            // code xB896 (tor-toong)
            16'h8960: data = 8'b00000000;
            16'h8961: data = 8'b00000000;
            16'h8962: data = 8'b00000000;
            16'h8963: data = 8'b00000000;
            16'h8964: data = 8'b00000000;
            16'h8965: data = 8'b01111000;
            16'h8966: data = 8'b11101100;
            16'h8967: data = 8'b01000110;
            16'h8968: data = 8'b11000110;
            16'h8969: data = 8'b11100110;
            16'h896A: data = 8'b10100110;
            16'h896B: data = 8'b11100110;
            16'h896C: data = 8'b00000000;
            16'h896D: data = 8'b00000000;
            16'h896E: data = 8'b00000000;
            16'h896F: data = 8'b00000000;
            
            // code xB897 (thor-tha-han)
            16'h8970: data = 8'b00000000;
            16'h8971: data = 8'b00000000;
            16'h8972: data = 8'b00000000;
            16'h8973: data = 8'b00000000;
            16'h8974: data = 8'b00000000;
            16'h8975: data = 8'b01000110;
            16'h8976: data = 8'b10100110;
            16'h8977: data = 8'b01101110;
            16'h8978: data = 8'b01111110;
            16'h8979: data = 8'b01110110;
            16'h897A: data = 8'b01100110;
            16'h897B: data = 8'b01100110;
            16'h897C: data = 8'b00000000;
            16'h897D: data = 8'b00000000;
            16'h897E: data = 8'b00000000;
            16'h897F: data = 8'b00000000;
            
            // code xB898 (tor-tong)
            16'h8980: data = 8'b00000000;
            16'h8981: data = 8'b00000000;
            16'h8982: data = 8'b00000000;
            16'h8983: data = 8'b00000000;
            16'h8984: data = 8'b00000000;
            16'h8985: data = 8'b01111110;
            16'h8986: data = 8'b11000000;
            16'h8987: data = 8'b11111100;
            16'h8988: data = 8'b00100110;
            16'h8989: data = 8'b01100110;
            16'h898A: data = 8'b01100110;
            16'h898B: data = 8'b01111100;
            16'h898C: data = 8'b00000000;
            16'h898D: data = 8'b00000000;
            16'h898E: data = 8'b00000000;
            16'h898F: data = 8'b00000000;
            
            // code xB899 (nor-nu)
            16'h8990: data = 8'b00000000;
            16'h8991: data = 8'b00000000;
            16'h8992: data = 8'b00000000;
            16'h8993: data = 8'b00000000;
            16'h8994: data = 8'b00000000;
            16'h8995: data = 8'b01000110;
            16'h8996: data = 8'b10100110;
            16'h8997: data = 8'b11100110;
            16'h8998: data = 8'b01100110;
            16'h8999: data = 8'b01001100;
            16'h899A: data = 8'b01111010;
            16'h899B: data = 8'b01100100;
            16'h899C: data = 8'b00000000;
            16'h899D: data = 8'b00000000;
            16'h899E: data = 8'b00000000;
            16'h899F: data = 8'b00000000;
            
            // code xB89A (bor-bai-mai)
            16'h89A0: data = 8'b00000000;
            16'h89A1: data = 8'b00000000;
            16'h89A2: data = 8'b00000000;
            16'h89A3: data = 8'b00000000;
            16'h89A4: data = 8'b00000000;
            16'h89A5: data = 8'b01000110;
            16'h89A6: data = 8'b10100110;
            16'h89A7: data = 8'b11100110;
            16'h89A8: data = 8'b01100110;
            16'h89A9: data = 8'b01100110;
            16'h89AA: data = 8'b01100110;
            16'h89AB: data = 8'b11111100;
            16'h89AC: data = 8'b00000000;
            16'h89AD: data = 8'b00000000;
            16'h89AE: data = 8'b00000000;
            16'h89AF: data = 8'b00000000;
            
            // code xB89B (por-pla)
            16'h89B0: data = 8'b00000000;
            16'h89B1: data = 8'b00000000;
            16'h89B2: data = 8'b00000110;
            16'h89B3: data = 8'b00000110;
            16'h89B4: data = 8'b00000110;
            16'h89B5: data = 8'b01000110;
            16'h89B6: data = 8'b10100110;
            16'h89B7: data = 8'b11100110;
            16'h89B8: data = 8'b01100110;
            16'h89B9: data = 8'b01100110;
            16'h89BA: data = 8'b01100110;
            16'h89BB: data = 8'b11111100;
            16'h89BC: data = 8'b00000000;
            16'h89BD: data = 8'b00000000;
            16'h89BE: data = 8'b00000000;
            16'h89BF: data = 8'b00000000;
            
            // code xB89C (phor-pueng)
            16'h89C0: data = 8'b00000000;
            16'h89C1: data = 8'b00000000;
            16'h89C2: data = 8'b00000000;
            16'h89C3: data = 8'b00000000;
            16'h89C4: data = 8'b00000000;
            16'h89C5: data = 8'b01000110;
            16'h89C6: data = 8'b10100110;
            16'h89C7: data = 8'b11000110;
            16'h89C8: data = 8'b11010110;
            16'h89C9: data = 8'b11111110;
            16'h89CA: data = 8'b11101110;
            16'h89CB: data = 8'b11100110;
            16'h89CC: data = 8'b00000000;
            16'h89CD: data = 8'b00000000;
            16'h89CE: data = 8'b00000000;
            16'h89CF: data = 8'b00000000;
            
            // code xB89D (phor-pueng)
            16'h89D0: data = 8'b00000000;
            16'h89D1: data = 8'b00000000;
            16'h89D2: data = 8'b00000000;
            16'h89D3: data = 8'b00000110;
            16'h89D4: data = 8'b00000110;
            16'h89D5: data = 8'b01000110;
            16'h89D6: data = 8'b10100110;
            16'h89D7: data = 8'b11000110;
            16'h89D8: data = 8'b11010110;
            16'h89D9: data = 8'b11111110;
            16'h89DA: data = 8'b11101110;
            16'h89DB: data = 8'b11100110;
            16'h89DC: data = 8'b00000000;
            16'h89DD: data = 8'b00000000;
            16'h89DE: data = 8'b00000000;
            16'h89DF: data = 8'b00000000;
            
            // code xB89E (por-phan)
            16'h89E0: data = 8'b00000000;
            16'h89E1: data = 8'b00000000;
            16'h89E2: data = 8'b00000000;
            16'h89E3: data = 8'b00000000;
            16'h89E4: data = 8'b00000000;
            16'h89E5: data = 8'b01000110;
            16'h89E6: data = 8'b10100110;
            16'h89E7: data = 8'b11100110;
            16'h89E8: data = 8'b01010110;
            16'h89E9: data = 8'b01111110;
            16'h89EA: data = 8'b01101110;
            16'h89EB: data = 8'b01100110;
            16'h89EC: data = 8'b00000000;
            16'h89ED: data = 8'b00000000;
            16'h89EE: data = 8'b00000000;
            16'h89EF: data = 8'b00000000;
            
            // code xB89F (for-fhan)
            16'h89F0: data = 8'b00000000;
            16'h89F1: data = 8'b00000000;
            16'h89F2: data = 8'b00000110;
            16'h89F3: data = 8'b00000110;
            16'h89F4: data = 8'b00000110;
            16'h89F5: data = 8'b01000110;
            16'h89F6: data = 8'b10100110;
            16'h89F7: data = 8'b11100110;
            16'h89F8: data = 8'b01010110;
            16'h89F9: data = 8'b01111110;
            16'h89FA: data = 8'b01101110;
            16'h89FB: data = 8'b01100110;
            16'h89FC: data = 8'b00000000;
            16'h89FD: data = 8'b00000000;
            16'h89FE: data = 8'b00000000;
            16'h89FF: data = 8'b00000000;
            
            16'h8976: data = 8'b00000000;	//
            16'h8977: data = 8'b00000000;	//
            16'h8978: data = 8'b00000000;	//
            16'h8979: data = 8'b00000000;	//
            16'h897A: data = 8'b00000000;	//
            16'h897B: data = 8'b00000000;	//
            16'h897C: data = 8'b00000000;	//
            16'h897D: data = 8'b00000000;	//
            16'h897E: data = 8'b00000000;	//
            16'h897F: data = 8'b00000000;	//
            
            // code xB898 (tor-tong)
            16'h8980: data = 8'b00000000;
            16'h8981: data = 8'b00000000;
            16'h8982: data = 8'b00000000;
            16'h8983: data = 8'b00000000;
            16'h8984: data = 8'b00000000;
            16'h8985: data = 8'b01111110;
            16'h8986: data = 8'b11000000;
            16'h8987: data = 8'b11111100;
            16'h8988: data = 8'b00100110;
            16'h8989: data = 8'b01100110;
            16'h898A: data = 8'b01100110;
            16'h898B: data = 8'b01111100;
            16'h898C: data = 8'b00000000;
            16'h898D: data = 8'b00000000;
            16'h898E: data = 8'b00000000;
            16'h898F: data = 8'b00000000;
            
            // code xB899 (nor-nu)
            16'h8990: data = 8'b00000000;
            16'h8991: data = 8'b00000000;
            16'h8992: data = 8'b00000000;
            16'h8993: data = 8'b00000000;
            16'h8994: data = 8'b00000000;
            16'h8995: data = 8'b01000110;
            16'h8996: data = 8'b10100110;
            16'h8997: data = 8'b11100110;
            16'h8998: data = 8'b01100110;
            16'h8999: data = 8'b01001100;
            16'h899A: data = 8'b01111010;
            16'h899B: data = 8'b01100100;
            16'h899C: data = 8'b00000000;
            16'h899D: data = 8'b00000000;
            16'h899E: data = 8'b00000000;
            16'h899F: data = 8'b00000000;
            
            // code xB89A (bor-bai-mai)
            16'h89A0: data = 8'b00000000;
            16'h89A1: data = 8'b00000000;
            16'h89A2: data = 8'b00000000;
            16'h89A3: data = 8'b00000000;
            16'h89A4: data = 8'b00000000;
            16'h89A5: data = 8'b01000110;
            16'h89A6: data = 8'b10100110;
            16'h89A7: data = 8'b11100110;
            16'h89A8: data = 8'b01100110;
            16'h89A9: data = 8'b01100110;
            16'h89AA: data = 8'b01100110;
            16'h89AB: data = 8'b11111100;
            16'h89AC: data = 8'b00000000;
            16'h89AD: data = 8'b00000000;
            16'h89AE: data = 8'b00000000;
            16'h89AF: data = 8'b00000000;
            
            // code xB89B (por-pla)
            16'h89B0: data = 8'b00000000;
            16'h89B1: data = 8'b00000000;
            16'h89B2: data = 8'b00000110;
            16'h89B3: data = 8'b00000110;
            16'h89B4: data = 8'b00000110;
            16'h89B5: data = 8'b01000110;
            16'h89B6: data = 8'b10100110;
            16'h89B7: data = 8'b11100110;
            16'h89B8: data = 8'b01100110;
            16'h89B9: data = 8'b01100110;
            16'h89BA: data = 8'b01100110;
            16'h89BB: data = 8'b11111100;
            16'h89BC: data = 8'b00000000;
            16'h89BD: data = 8'b00000000;
            16'h89BE: data = 8'b00000000;
            16'h89BF: data = 8'b00000000;
            
            // code xB89C (t28)
            16'h89C0: data = 8'b00000000;	//
            16'h89C1: data = 8'b00000000;	//
            16'h89C2: data = 8'b00000000;	//
            16'h89C3: data = 8'b00000000;	//
            16'h89C4: data = 8'b00000000;	//
            16'h89C5: data = 8'b00000000;	//
            16'h89C6: data = 8'b00000000;	//
            16'h89C7: data = 8'b00000000;	//
            16'h89C8: data = 8'b00000000;	//
            16'h89C9: data = 8'b00000000;	//
            16'h89CA: data = 8'b00000000;	//
            16'h89CB: data = 8'b00000000;	//
            16'h89CC: data = 8'b00000000;	//
            16'h89CD: data = 8'b00000000;	//
            16'h89CE: data = 8'b00000000;	//
            16'h89CF: data = 8'b00000000;	//
            
            // code xB89D (t29)
            16'h89D0: data = 8'b00000000;	//
            16'h89D1: data = 8'b00000000;	//
            16'h89D2: data = 8'b00000000;	//
            16'h89D3: data = 8'b00000000;	//
            16'h89D4: data = 8'b00000000;	//
            16'h89D5: data = 8'b00000000;	//
            16'h89D6: data = 8'b00000000;	//
            16'h89D7: data = 8'b00000000;	//
            16'h89D8: data = 8'b00000000;	//
            16'h89D9: data = 8'b00000000;	//
            16'h89DA: data = 8'b00000000;	//
            16'h89DB: data = 8'b00000000;	//
            16'h89DC: data = 8'b00000000;	//
            16'h89DD: data = 8'b00000000;	//
            16'h89DE: data = 8'b00000000;	//
            16'h89DF: data = 8'b00000000;	//
            
            // code xB89E (t30)
            16'h89E0: data = 8'b00000000;	//
            16'h89E1: data = 8'b00000000;	//
            16'h89E2: data = 8'b00000000;	//
            16'h89E3: data = 8'b00000000;	//
            16'h89E4: data = 8'b00000000;	//
            16'h89E5: data = 8'b00000000;	//
            16'h89E6: data = 8'b00000000;	//
            16'h89E7: data = 8'b00000000;	//
            16'h89E8: data = 8'b00000000;	//
            16'h89E9: data = 8'b00000000;	//
            16'h89EA: data = 8'b00000000;	//
            16'h89EB: data = 8'b00000000;	//
            16'h89EC: data = 8'b00000000;	//
            16'h89ED: data = 8'b00000000;	//
            16'h89EE: data = 8'b00000000;	//
            16'h89EF: data = 8'b00000000;	//
            
            // code xB89F (t31)
            16'h89F0: data = 8'b00000000;	//
            16'h89F1: data = 8'b00000000;	//
            16'h89F2: data = 8'b00000000;	//
            16'h89F3: data = 8'b00000000;	//
            16'h89F4: data = 8'b00000000;	//
            16'h89F5: data = 8'b00000000;	//
            16'h89F6: data = 8'b00000000;	//
            16'h89F7: data = 8'b00000000;	//
            16'h89F8: data = 8'b00000000;	//
            16'h89F9: data = 8'b00000000;	//
            16'h89FA: data = 8'b00000000;	//
            16'h89FB: data = 8'b00000000;	//
            16'h89FC: data = 8'b00000000;	//
            16'h89FD: data = 8'b00000000;	//
            16'h89FE: data = 8'b00000000;	//
            16'h89FF: data = 8'b00000000;	//
            
            // code xB8A0 (por-sum-pao)
            16'h8A00: data = 8'b00000000;
            16'h8A01: data = 8'b00000000;
            16'h8A02: data = 8'b00000000;
            16'h8A03: data = 8'b00000000;
            16'h8A04: data = 8'b00000000;
            16'h8A05: data = 8'b00111100;
            16'h8A06: data = 8'b01111110;
            16'h8A07: data = 8'b11100110;
            16'h8A08: data = 8'b00100110;
            16'h8A09: data = 8'b01100110;
            16'h8A0A: data = 8'b10100110;
            16'h8A0B: data = 8'b01100110;
            16'h8A0C: data = 8'b00000000;
            16'h8A0D: data = 8'b00000000;
            16'h8A0E: data = 8'b00000000;
            16'h8A0F: data = 8'b00000000;
            
            // code xB8A1 (mor-mar)
            16'h8A10: data = 8'b00000000;
            16'h8A11: data = 8'b00000000;
            16'h8A12: data = 8'b00000000;
            16'h8A13: data = 8'b00000000;
            16'h8A14: data = 8'b00000000;
            16'h8A15: data = 8'b01000110;
            16'h8A16: data = 8'b10100110;
            16'h8A17: data = 8'b01100110;
            16'h8A18: data = 8'b01100110;
            16'h8A19: data = 8'b01110110;
            16'h8A1A: data = 8'b10101110;
            16'h8A1B: data = 8'b01100110;
            16'h8A1C: data = 8'b00000000;
            16'h8A1D: data = 8'b00000000;
            16'h8A1E: data = 8'b00000000;
            16'h8A1F: data = 8'b00000000;
            
            // code xB8A2 (yor-yak)
            16'h8A20: data = 8'b00000000;
            16'h8A21: data = 8'b00000000;
            16'h8A22: data = 8'b00000000;
            16'h8A23: data = 8'b00000000;
            16'h8A24: data = 8'b00000000;
            16'h8A25: data = 8'b01000110;
            16'h8A26: data = 8'b10100110;
            16'h8A27: data = 8'b11000110;
            16'h8A28: data = 8'b01100110;
            16'h8A29: data = 8'b11000110;
            16'h8A2A: data = 8'b11101110;
            16'h8A2B: data = 8'b01111100;
            16'h8A2C: data = 8'b00000000;
            16'h8A2D: data = 8'b00000000;
            16'h8A2E: data = 8'b00000000;
            16'h8A2F: data = 8'b00000000;
            
            // code xB8A3 (ror-rue)
            16'h8A30: data = 8'b00000000;
            16'h8A31: data = 8'b00000000;
            16'h8A32: data = 8'b00000000;
            16'h8A33: data = 8'b00000000;
            16'h8A34: data = 8'b00000000;
            16'h8A35: data = 8'b01111110;
            16'h8A36: data = 8'b11000000;
            16'h8A37: data = 8'b11110000;
            16'h8A38: data = 8'b00111000;
            16'h8A39: data = 8'b00011000;
            16'h8A3A: data = 8'b00101000;
            16'h8A3B: data = 8'b00011000;
            16'h8A3C: data = 8'b00000000;
            16'h8A3D: data = 8'b00000000;
            16'h8A3E: data = 8'b00000000;
            16'h8A3F: data = 8'b00000000;
            
            // code xB8A4 (ror-rue-1)
            16'h8A40: data = 8'b00000000;
            16'h8A41: data = 8'b00000000;
            16'h8A42: data = 8'b00000000;
            16'h8A43: data = 8'b00000000;
            16'h8A44: data = 8'b00000000;
            16'h8A45: data = 8'b01111100;
            16'h8A46: data = 8'b11001100;
            16'h8A47: data = 8'b01000110;
            16'h8A48: data = 8'b11000110;
            16'h8A49: data = 8'b11000110;
            16'h8A4A: data = 8'b10100110;
            16'h8A4B: data = 8'b01100110;
            16'h8A4C: data = 8'b00000110;
            16'h8A4D: data = 8'b00000110;
            16'h8A4E: data = 8'b00000110;
            16'h8A4F: data = 8'b00000000;
            
            // code xB8A5 (lor-ling)
            16'h8A50: data = 8'b00000000;
            16'h8A51: data = 8'b00000000;
            16'h8A52: data = 8'b00000000;
            16'h8A53: data = 8'b00000000;
            16'h8A54: data = 8'b00000000;
            16'h8A55: data = 8'b01111100;
            16'h8A56: data = 8'b11001100;
            16'h8A57: data = 8'b11000110;
            16'h8A58: data = 8'b00110110;
            16'h8A59: data = 8'b01111110;
            16'h8A5A: data = 8'b10101110;
            16'h8A5B: data = 8'b01100110;
            16'h8A5C: data = 8'b00000000;
            16'h8A5D: data = 8'b00000000;
            16'h8A5E: data = 8'b00000000;
            16'h8A5F: data = 8'b00000000;
            
            // code xB8A6 (ror-long)
            16'h8A60: data = 8'b00000000;
            16'h8A61: data = 8'b00000000;
            16'h8A62: data = 8'b00000000;
            16'h8A63: data = 8'b00000000;
            16'h8A64: data = 8'b00000000;
            16'h8A65: data = 8'b01111100;
            16'h8A66: data = 8'b11001100;
            16'h8A67: data = 8'b11000110;
            16'h8A68: data = 8'b01100110;
            16'h8A69: data = 8'b01100110;
            16'h8A6A: data = 8'b10100110;
            16'h8A6B: data = 8'b01100110;
            16'h8A6C: data = 8'b00000110;
            16'h8A6D: data = 8'b00000110;
            16'h8A6E: data = 8'b00000110;
            16'h8A6F: data = 8'b00000000;
            
            // code xB8A7 (vor-van)
            16'h8A70: data = 8'b00000000;
            16'h8A71: data = 8'b00000000;
            16'h8A72: data = 8'b00000000;
            16'h8A73: data = 8'b00000000;
            16'h8A74: data = 8'b00000000;
            16'h8A75: data = 8'b00111100;
            16'h8A76: data = 8'b01101110;
            16'h8A77: data = 8'b11000110;
            16'h8A78: data = 8'b00000110;
            16'h8A79: data = 8'b00001110;
            16'h8A7A: data = 8'b00010110;
            16'h8A7B: data = 8'b00011100;
            16'h8A7C: data = 8'b00000000;
            16'h8A7D: data = 8'b00000000;
            16'h8A7E: data = 8'b00000000;
            16'h8A7F: data = 8'b00000000;
            
            // code xB8A8 (sor-1)
            16'h8A80: data = 8'b00000000;
            16'h8A81: data = 8'b00000000;
            16'h8A82: data = 8'b00000000;
            16'h8A83: data = 8'b00000010;
            16'h8A84: data = 8'b00000110;
            16'h8A85: data = 8'b00111100;
            16'h8A86: data = 8'b01101100;
            16'h8A87: data = 8'b11000110;
            16'h8A88: data = 8'b11010110;
            16'h8A89: data = 8'b11101110;
            16'h8A8A: data = 8'b11110110;
            16'h8A8B: data = 8'b11000110;
            16'h8A8C: data = 8'b00000000;
            16'h8A8D: data = 8'b00000000;
            16'h8A8E: data = 8'b00000000;
            16'h8A8F: data = 8'b00000000;
            
            // code xB8A9 (sor-2)
            16'h8A90: data = 8'b00000000;
            16'h8A91: data = 8'b00000000;
            16'h8A92: data = 8'b00000000;
            16'h8A93: data = 8'b00000000;
            16'h8A94: data = 8'b00000000;
            16'h8A95: data = 8'b01000110;
            16'h8A96: data = 8'b10100110;
            16'h8A97: data = 8'b01101110;
            16'h8A98: data = 8'b01010111;
            16'h8A99: data = 8'b01101111;
            16'h8A9A: data = 8'b01100110;
            16'h8A9B: data = 8'b11111110;
            16'h8A9C: data = 8'b00000000;
            16'h8A9D: data = 8'b00000000;
            16'h8A9E: data = 8'b00000000;
            16'h8A9F: data = 8'b00000000;
            
            // code xB8AA (sor-3)
            16'h8AA0: data = 8'b00000000;
            16'h8AA1: data = 8'b00000000;
            16'h8AA2: data = 8'b00000000;
            16'h8AA3: data = 8'b00000010;
            16'h8AA4: data = 8'b00000010;
            16'h8AA5: data = 8'b00111100;
            16'h8AA6: data = 8'b01101100;
            16'h8AA7: data = 8'b11000110;
            16'h8AA8: data = 8'b00000110;
            16'h8AA9: data = 8'b01111110;
            16'h8AAA: data = 8'b10101110;
            16'h8AAB: data = 8'b01100110;
            16'h8AAC: data = 8'b00000000;
            16'h8AAD: data = 8'b00000000;
            16'h8AAE: data = 8'b00000000;
            16'h8AAF: data = 8'b00000000;
            
            // code xB8AB (hor-heep)
            16'h8AB0: data = 8'b00000000;
            16'h8AB1: data = 8'b00000000;
            16'h8AB2: data = 8'b00000000;
            16'h8AB3: data = 8'b00000000;
            16'h8AB4: data = 8'b00000000;
            16'h8AB5: data = 8'b01100110;
            16'h8AB6: data = 8'b10101010;
            16'h8AB7: data = 8'b01101100;
            16'h8AB8: data = 8'b00110110;
            16'h8AB9: data = 8'b01100110;
            16'h8ABA: data = 8'b01100110;
            16'h8ABB: data = 8'b01100110;
            16'h8ABC: data = 8'b00000000;
            16'h8ABD: data = 8'b00000000;
            16'h8ABE: data = 8'b00000000;
            16'h8ABF: data = 8'b00000000;
            
            // code xB8AC (chula)
            16'h8AC0: data = 8'b00000000;
            16'h8AC1: data = 8'b00000000;
            16'h8AC2: data = 8'b00000001;
            16'h8AC3: data = 8'b00000111;
            16'h8AC4: data = 8'b00001010;
            16'h8AC5: data = 8'b01000110;
            16'h8AC6: data = 8'b10100110;
            16'h8AC7: data = 8'b01100110;
            16'h8AC8: data = 8'b01010110;
            16'h8AC9: data = 8'b01111110;
            16'h8ACA: data = 8'b01101110;
            16'h8ACB: data = 8'b01000110;
            16'h8ACC: data = 8'b00000000;
            16'h8ACD: data = 8'b00000000;
            16'h8ACE: data = 8'b00000000;
            16'h8ACF: data = 8'b00000000;
            
            // code xB8AD (oor)
            16'h8AD0: data = 8'b00000000;
            16'h8AD1: data = 8'b00000000;
            16'h8AD2: data = 8'b00000000;
            16'h8AD3: data = 8'b00000000;
            16'h8AD4: data = 8'b00000000;
            16'h8AD5: data = 8'b01111000;
            16'h8AD6: data = 8'b11001100;
            16'h8AD7: data = 8'b00000110;
            16'h8AD8: data = 8'b11100110;
            16'h8AD9: data = 8'b10100110;
            16'h8ADA: data = 8'b11000110;
            16'h8ADB: data = 8'b11111110;
            16'h8ADC: data = 8'b00000000;
            16'h8ADD: data = 8'b00000000;
            16'h8ADE: data = 8'b00000000;
            16'h8ADF: data = 8'b00000000;
            
            // code xB8AE (hor-nok-hoog)
            16'h8AE0: data = 8'b00000000;
            16'h8AE1: data = 8'b00000000;
            16'h8AE2: data = 8'b00000000;
            16'h8AE3: data = 8'b00000010;
            16'h8AE4: data = 8'b00000110;
            16'h8AE5: data = 8'b01111100;
            16'h8AE6: data = 8'b11001100;
            16'h8AE7: data = 8'b00000110;
            16'h8AE8: data = 8'b11100110;
            16'h8AE9: data = 8'b10100110;
            16'h8AEA: data = 8'b11000110;
            16'h8AEB: data = 8'b11111110;
            16'h8AEC: data = 8'b00000000;
            16'h8AED: data = 8'b00000000;
            16'h8AEE: data = 8'b00000000;
            16'h8AEF: data = 8'b00000000;
            
            // code xB8AF (pai-yarn)
            16'h8AF0: data = 8'b00000000;
            16'h8AF1: data = 8'b00000000;
            16'h8AF2: data = 8'b00000000;
            16'h8AF3: data = 8'b00000000;
            16'h8AF4: data = 8'b00000000;
            16'h8AF5: data = 8'b01100110;
            16'h8AF6: data = 8'b10101110;
            16'h8AF7: data = 8'b01111110;
            16'h8AF8: data = 8'b00000110;
            16'h8AF9: data = 8'b00000110;
            16'h8AFA: data = 8'b00000110;
            16'h8AFB: data = 8'b00001100;
            16'h8AFC: data = 8'b00000000;
            16'h8AFD: data = 8'b00000000;
            16'h8AFE: data = 8'b00000000;
            16'h8AFF: data = 8'b00000000;
            
            // code xB8B0 (a)
            16'h8B00: data = 8'b00000000;
            16'h8B01: data = 8'b00000000;
            16'h8B02: data = 8'b00000000;
            16'h8B03: data = 8'b00000000;
            16'h8B04: data = 8'b00000000;
            16'h8B05: data = 8'b01000010;
            16'h8B06: data = 8'b10100110;
            16'h8B07: data = 8'b11111100;
            16'h8B08: data = 8'b01000010;
            16'h8B09: data = 8'b10100110;
            16'h8B0A: data = 8'b11111100;
            16'h8B0B: data = 8'b00000000;
            16'h8B0C: data = 8'b00000000;
            16'h8B0D: data = 8'b00000000;
            16'h8B0E: data = 8'b00000000;
            16'h8B0F: data = 8'b00000000;
            
            // code xB8B1 (a-2)
            16'h8B10: data = 8'b00000000;
            16'h8B11: data = 8'b00100010;
            16'h8B12: data = 8'b01010110;
            16'h8B13: data = 8'b01111100;
            16'h8B14: data = 8'b00000000;
            16'h8B15: data = 8'b00000000;
            16'h8B16: data = 8'b00000000;
            16'h8B17: data = 8'b00000000;
            16'h8B18: data = 8'b00000000;
            16'h8B19: data = 8'b00000000;
            16'h8B1A: data = 8'b00000000;
            16'h8B1B: data = 8'b00000000;
            16'h8B1C: data = 8'b00000000;
            16'h8B1D: data = 8'b00000000;
            16'h8B1E: data = 8'b00000000;
            16'h8B1F: data = 8'b00000000;
            
            // code xB8B2 (ar)
            16'h8B20: data = 8'b00000000;
            16'h8B21: data = 8'b00000000;
            16'h8B22: data = 8'b00000000;
            16'h8B23: data = 8'b00000000;
            16'h8B24: data = 8'b00000000;
            16'h8B25: data = 8'b00111000;
            16'h8B26: data = 8'b01111100;
            16'h8B27: data = 8'b01001110;
            16'h8B28: data = 8'b00000110;
            16'h8B29: data = 8'b00000110;
            16'h8B2A: data = 8'b00000110;
            16'h8B2B: data = 8'b00000110;
            16'h8B2C: data = 8'b00000000;
            16'h8B2D: data = 8'b00000000;
            16'h8B2E: data = 8'b00000000;
            16'h8B2F: data = 8'b00000000;
            
            // code xB8B3 (aum)
            16'h8B30: data = 8'b00000000;
            16'h8B31: data = 8'b01000000;
            16'h8B32: data = 8'b10100000;
            16'h8B33: data = 8'b01000000;
            16'h8B34: data = 8'b00000000;
            16'h8B35: data = 8'b00111000;
            16'h8B36: data = 8'b01111100;
            16'h8B37: data = 8'b01001110;
            16'h8B38: data = 8'b00000110;
            16'h8B39: data = 8'b00000110;
            16'h8B3A: data = 8'b00000110;
            16'h8B3B: data = 8'b00000110;
            16'h8B3C: data = 8'b00000000;
            16'h8B3D: data = 8'b00000000;
            16'h8B3E: data = 8'b00000000;
            16'h8B3F: data = 8'b00000000;
            
            // code xB8B4 (ei)
            16'h8B40: data = 8'b00000000;
            16'h8B41: data = 8'b00110000;
            16'h8B42: data = 8'b01001000;
            16'h8B43: data = 8'b01111000;
            16'h8B44: data = 8'b00000000;
            16'h8B45: data = 8'b00000000;
            16'h8B46: data = 8'b00000000;
            16'h8B47: data = 8'b00000000;
            16'h8B48: data = 8'b00000000;
            16'h8B49: data = 8'b00000000;
            16'h8B4A: data = 8'b00000000;
            16'h8B4B: data = 8'b00000000;
            16'h8B4C: data = 8'b00000000;
            16'h8B4D: data = 8'b00000000;
            16'h8B4E: data = 8'b00000000;
            16'h8B4F: data = 8'b00000000;
            
            // code xB8B5 (ee)
            16'h8B50: data = 8'b00000000;
            16'h8B51: data = 8'b00110100;
            16'h8B52: data = 8'b01001100;
            16'h8B53: data = 8'b01111100;
            16'h8B54: data = 8'b00000000;
            16'h8B55: data = 8'b00000000;
            16'h8B56: data = 8'b00000000;
            16'h8B57: data = 8'b00000000;
            16'h8B58: data = 8'b00000000;
            16'h8B59: data = 8'b00000000;
            16'h8B5A: data = 8'b00000000;
            16'h8B5B: data = 8'b00000000;
            16'h8B5C: data = 8'b00000000;
            16'h8B5D: data = 8'b00000000;
            16'h8B5E: data = 8'b00000000;
            16'h8B5F: data = 8'b00000000;
            
            // code xB8B6 (ue)
            16'h8B60: data = 8'b00000000;
            16'h8B61: data = 8'b00110100;
            16'h8B62: data = 8'b01001010;
            16'h8B63: data = 8'b01111100;
            16'h8B64: data = 8'b00000000;
            16'h8B65: data = 8'b00000000;
            16'h8B66: data = 8'b00000000;
            16'h8B67: data = 8'b00000000;
            16'h8B68: data = 8'b00000000;
            16'h8B69: data = 8'b00000000;
            16'h8B6A: data = 8'b00000000;
            16'h8B6B: data = 8'b00000000;
            16'h8B6C: data = 8'b00000000;
            16'h8B6D: data = 8'b00000000;
            16'h8B6E: data = 8'b00000000;
            16'h8B6F: data = 8'b00000000;
            
            // code xB8B7 (uee)
            16'h8B70: data = 8'b00000000;
            16'h8B71: data = 8'b00101010;
            16'h8B72: data = 8'b01011010;
            16'h8B73: data = 8'b01111110;
            16'h8B74: data = 8'b00000000;
            16'h8B75: data = 8'b00000000;
            16'h8B76: data = 8'b00000000;
            16'h8B77: data = 8'b00000000;
            16'h8B78: data = 8'b00000000;
            16'h8B79: data = 8'b00000000;
            16'h8B7A: data = 8'b00000000;
            16'h8B7B: data = 8'b00000000;
            16'h8B7C: data = 8'b00000000;
            16'h8B7D: data = 8'b00000000;
            16'h8B7E: data = 8'b00000000;
            16'h8B7F: data = 8'b00000000;
            
            // code xB8B8 (u)
            16'h8B80: data = 8'b00000000;
            16'h8B81: data = 8'b00000000;
            16'h8B82: data = 8'b00000000;
            16'h8B83: data = 8'b00000000;
            16'h8B84: data = 8'b00000000;
            16'h8B85: data = 8'b00000000;
            16'h8B86: data = 8'b00000000;
            16'h8B87: data = 8'b00000000;
            16'h8B88: data = 8'b00000000;
            16'h8B89: data = 8'b00000000;
            16'h8B8A: data = 8'b00000000;
            16'h8B8B: data = 8'b00000000;
            16'h8B8C: data = 8'b00010000;
            16'h8B8D: data = 8'b00101000;
            16'h8B8E: data = 8'b00011000;
            16'h8B8F: data = 8'b00001000;
            
            // code xB8B9 (uu)
            16'h8B90: data = 8'b00000000;
            16'h8B91: data = 8'b00000000;
            16'h8B92: data = 8'b00000000;
            16'h8B93: data = 8'b00000000;
            16'h8B94: data = 8'b00000000;
            16'h8B95: data = 8'b00000000;
            16'h8B96: data = 8'b00000000;
            16'h8B97: data = 8'b00000000;
            16'h8B98: data = 8'b00000000;
            16'h8B99: data = 8'b00000000;
            16'h8B9A: data = 8'b00000000;
            16'h8B9B: data = 8'b00000000;
            16'h8B9C: data = 8'b00110100;
            16'h8B9D: data = 8'b01010100;
            16'h8B9E: data = 8'b00110100;
            16'h8B9F: data = 8'b00011000;
            
            // code xB8BA (phinthu)
            16'h8BA0: data = 8'b00000000;
            16'h8BA1: data = 8'b00000000;
            16'h8BA2: data = 8'b00000000;
            16'h8BA3: data = 8'b00000000;
            16'h8BA4: data = 8'b00000000;
            16'h8BA5: data = 8'b00000000;
            16'h8BA6: data = 8'b00000000;
            16'h8BA7: data = 8'b00000000;
            16'h8BA8: data = 8'b00000000;
            16'h8BA9: data = 8'b00000000;
            16'h8BAA: data = 8'b00000000;
            16'h8BAB: data = 8'b00000000;
            16'h8BAC: data = 8'b00000000;
            16'h8BAD: data = 8'b00000110;
            16'h8BAE: data = 8'b00000110;
            16'h8BAF: data = 8'b00000000;
            
            // code xB83F (baht)
            16'h83F0: data = 8'b00000000;
            16'h83F1: data = 8'b00000000;
            16'h83F2: data = 8'b00000000;
            16'h83F3: data = 8'b00000000;
            16'h83F4: data = 8'b00100000;
            16'h83F5: data = 8'b11111000;
            16'h83F6: data = 8'b10101100;
            16'h83F7: data = 8'b10100110;
            16'h83F8: data = 8'b10101100;
            16'h83F9: data = 8'b10101100;
            16'h83FA: data = 8'b10100110;
            16'h83FB: data = 8'b10101100;
            16'h83FC: data = 8'b11111000;
            16'h83FD: data = 8'b00100000;
            16'h83FE: data = 8'b00000000;
            16'h83FF: data = 8'b00000000;
            
            // code xB980 (e)
            16'h9800: data = 8'b00000000;
            16'h9801: data = 8'b00000000;
            16'h9802: data = 8'b00000000;
            16'h9803: data = 8'b00000000;
            16'h9804: data = 8'b00000000;
            16'h9805: data = 8'b00100000;
            16'h9806: data = 8'b00100000;
            16'h9807: data = 8'b00100000;
            16'h9808: data = 8'b00100000;
            16'h9809: data = 8'b00110000;
            16'h980A: data = 8'b00101000;
            16'h980B: data = 8'b00010000;
            16'h980C: data = 8'b00000000;
            16'h980D: data = 8'b00000000;
            16'h980E: data = 8'b00000000;
            16'h980F: data = 8'b00000000;
            
            // code xB981 (ae)
            16'h9810: data = 8'b00000000;
            16'h9811: data = 8'b00000000;
            16'h9812: data = 8'b00000000;
            16'h9813: data = 8'b00000000;
            16'h9814: data = 8'b00000000;
            16'h9815: data = 8'b10001000;
            16'h9816: data = 8'b10001000;
            16'h9817: data = 8'b10001000;
            16'h9818: data = 8'b10001000;
            16'h9819: data = 8'b11001100;
            16'h981A: data = 8'b10101010;
            16'h981B: data = 8'b01000100;
            16'h981C: data = 8'b00000000;
            16'h981D: data = 8'b00000000;
            16'h981E: data = 8'b00000000;
            16'h981F: data = 8'b00000000;
            
            // code xB982 (o)
            16'h9820: data = 8'b00000000;
            16'h9821: data = 8'b00000000;
            16'h9822: data = 8'b01001110;
            16'h9823: data = 8'b10111000;
            16'h9824: data = 8'b11000000;
            16'h9825: data = 8'b01100000;
            16'h9826: data = 8'b00100000;
            16'h9827: data = 8'b00100000;
            16'h9828: data = 8'b00100000;
            16'h9829: data = 8'b00110000;
            16'h982A: data = 8'b00101000;
            16'h982B: data = 8'b00010000;
            16'h982C: data = 8'b00000000;
            16'h982D: data = 8'b00000000;
            16'h982E: data = 8'b00000000;
            16'h982F: data = 8'b00000000;
            
            // code xB983 (ai)
            16'h9830: data = 8'b00000000;
            16'h9831: data = 8'b00000000;
            16'h9832: data = 8'b00110000;
            16'h9833: data = 8'b01001000;
            16'h9834: data = 8'b10101000;
            16'h9835: data = 8'b01001000;
            16'h9836: data = 8'b00001000;
            16'h9837: data = 8'b00001000;
            16'h9838: data = 8'b00001000;
            16'h9839: data = 8'b00001100;
            16'h983A: data = 8'b00001010;
            16'h983B: data = 8'b00000100;
            16'h983C: data = 8'b00000000;
            16'h983D: data = 8'b00000000;
            16'h983E: data = 8'b00000000;
            16'h983F: data = 8'b00000000;
            
            // code xB984 (ai-lai)
            16'h9840: data = 8'b00000000;
            16'h9841: data = 8'b00000000;
            16'h9842: data = 8'b10010000;
            16'h9843: data = 8'b10101000;
            16'h9844: data = 8'b01001000;
            16'h9845: data = 8'b00001000;
            16'h9846: data = 8'b00001000;
            16'h9847: data = 8'b00001000;
            16'h9848: data = 8'b00001000;
            16'h9849: data = 8'b00001100;
            16'h984A: data = 8'b00001010;
            16'h984B: data = 8'b00000100;
            16'h984C: data = 8'b00000000;
            16'h984D: data = 8'b00000000;
            16'h984E: data = 8'b00000000;
            16'h984F: data = 8'b00000000;
            
            // code xB985 (ar-long)
            16'h9850: data = 8'b00000000;
            16'h9851: data = 8'b00000000;
            16'h9852: data = 8'b00000000;
            16'h9853: data = 8'b00000000;
            16'h9854: data = 8'b00000000;
            16'h9855: data = 8'b00111100;
            16'h9856: data = 8'b01100110;
            16'h9857: data = 8'b00000110;
            16'h9858: data = 8'b00000110;
            16'h9859: data = 8'b00000110;
            16'h985A: data = 8'b00000110;
            16'h985B: data = 8'b00000110;
            16'h985C: data = 8'b00000110;
            16'h985D: data = 8'b00000110;
            16'h985E: data = 8'b00000000;
            16'h985F: data = 8'b00000000;
            
            // code xB986 (maiyamok)
            16'h9860: data = 8'b00000000;
            16'h9861: data = 8'b00000000;
            16'h9862: data = 8'b00000000;
            16'h9863: data = 8'b00000000;
            16'h9864: data = 8'b00000000;
            16'h9865: data = 8'b00000000;
            16'h9866: data = 8'b00000000;
            16'h9867: data = 8'b01011000;
            16'h9868: data = 8'b10101100;
            16'h9869: data = 8'b10000110;
            16'h986A: data = 8'b01000110;
            16'h986B: data = 8'b00000110;
            16'h986C: data = 8'b00000110;
            16'h986D: data = 8'b00000110;
            16'h986E: data = 8'b00001100;
            16'h986F: data = 8'b00000000;
            
            // code xB987 (maitaikhu)
            16'h9870: data = 8'b00000100;
            16'h9871: data = 8'b00101100;
            16'h9872: data = 8'b01010100;
            16'h9873: data = 8'b00101000;
            16'h9874: data = 8'b00000000;
            16'h9875: data = 8'b00000000;
            16'h9876: data = 8'b00000000;
            16'h9877: data = 8'b00000000;
            16'h9878: data = 8'b00000000;
            16'h9879: data = 8'b00000000;
            16'h987A: data = 8'b00000000;
            16'h987B: data = 8'b00000000;
            16'h987C: data = 8'b00000000;
            16'h987D: data = 8'b00000000;
            16'h987E: data = 8'b00000000;
            16'h987F: data = 8'b00000000;
            
            // code xB988 (mai-ek)
            16'h9880: data = 8'b00000000;
            16'h9881: data = 8'b00000010;
            16'h9882: data = 8'b00000010;
            16'h9883: data = 8'b00000010;
            16'h9884: data = 8'b00000000;
            16'h9885: data = 8'b00000000;
            16'h9886: data = 8'b00000000;
            16'h9887: data = 8'b00000000;
            16'h9888: data = 8'b00000000;
            16'h9889: data = 8'b00000000;
            16'h988A: data = 8'b00000000;
            16'h988B: data = 8'b00000000;
            16'h988C: data = 8'b00000000;
            16'h988D: data = 8'b00000000;
            16'h988E: data = 8'b00000000;
            16'h988F: data = 8'b00000000;
            
            // code xB989 (mai-tho)
            16'h9890: data = 8'b00000000;
            16'h9891: data = 8'b00000010;
            16'h9892: data = 8'b00010110;
            16'h9893: data = 8'b00011100;
            16'h9894: data = 8'b00000000;
            16'h9895: data = 8'b00000000;
            16'h9896: data = 8'b00000000;
            16'h9897: data = 8'b00000000;
            16'h9898: data = 8'b00000000;
            16'h9899: data = 8'b00000000;
            16'h989A: data = 8'b00000000;
            16'h989B: data = 8'b00000000;
            16'h989C: data = 8'b00000000;
            16'h989D: data = 8'b00000000;
            16'h989E: data = 8'b00000000;
            16'h989F: data = 8'b00000000;
            
            // code xB98A (mai-tri)
            16'h98A0: data = 8'b00000010;
            16'h98A1: data = 8'b01010110;
            16'h98A2: data = 8'b10101110;
            16'h98A3: data = 8'b01001000;
            16'h98A4: data = 8'b00000000;
            16'h98A5: data = 8'b00000000;
            16'h98A6: data = 8'b00000000;
            16'h98A7: data = 8'b00000000;
            16'h98A8: data = 8'b00000000;
            16'h98A9: data = 8'b00000000;
            16'h98AA: data = 8'b00000000;
            16'h98AB: data = 8'b00000000;
            16'h98AC: data = 8'b00000000;
            16'h98AD: data = 8'b00000000;
            16'h98AE: data = 8'b00000000;
            16'h98AF: data = 8'b00000000;
            
            // code xB98B (mai-chattawa)
            16'h98B0: data = 8'b00000000;
            16'h98B1: data = 8'b00000100;
            16'h98B2: data = 8'b00001110;
            16'h98B3: data = 8'b00000100;
            16'h98B4: data = 8'b00000000;
            16'h98B5: data = 8'b00000000;
            16'h98B6: data = 8'b00000000;
            16'h98B7: data = 8'b00000000;
            16'h98B8: data = 8'b00000000;
            16'h98B9: data = 8'b00000000;
            16'h98BA: data = 8'b00000000;
            16'h98BB: data = 8'b00000000;
            16'h98BC: data = 8'b00000000;
            16'h98BD: data = 8'b00000000;
            16'h98BE: data = 8'b00000000;
            16'h98BF: data = 8'b00000000;
            
            // code xB98C (thanthakhat)
            16'h98C0: data = 8'b00000010;
            16'h98C1: data = 8'b00011110;
            16'h98C2: data = 8'b00101000;
            16'h98C3: data = 8'b00010000;
            16'h98C4: data = 8'b00000000;
            16'h98C5: data = 8'b00000000;
            16'h98C6: data = 8'b00000000;
            16'h98C7: data = 8'b00000000;
            16'h98C8: data = 8'b00000000;
            16'h98C9: data = 8'b00000000;
            16'h98CA: data = 8'b00000000;
            16'h98CB: data = 8'b00000000;
            16'h98CC: data = 8'b00000000;
            16'h98CD: data = 8'b00000000;
            16'h98CE: data = 8'b00000000;
            16'h98CF: data = 8'b00000000;
            // code x990 (0-TH)
            16'h9900: data = 8'b00000000;
            16'h9901: data = 8'b00000000;
            16'h9902: data = 8'b00000000;
            16'h9903: data = 8'b00111000;
            16'h9904: data = 8'b01111100;
            16'h9905: data = 8'b01000100;
            16'h9906: data = 8'b10000010;
            16'h9907: data = 8'b10000010;
            16'h9908: data = 8'b10000010;
            16'h9909: data = 8'b11000110;
            16'h990A: data = 8'b01111100;
            16'h990B: data = 8'b00111000;
            16'h990C: data = 8'b00000000;
            16'h990D: data = 8'b00000000;
            16'h990E: data = 8'b00000000;
            16'h990F: data = 8'b00000000;
            // code x991 (1-TH)
            16'h9910: data = 8'b00000000;
            16'h9911: data = 8'b00000000;
            16'h9912: data = 8'b00000000;
            16'h9913: data = 8'b00111000;
            16'h9914: data = 8'b01111100;
            16'h9915: data = 8'b01000100;
            16'h9916: data = 8'b10000010;
            16'h9917: data = 8'b10111010;
            16'h9918: data = 8'b10101010;
            16'h9919: data = 8'b01110010;
            16'h991A: data = 8'b00000110;
            16'h991B: data = 8'b00111100;
            16'h991C: data = 8'b00000000;
            16'h991D: data = 8'b00000000;
            16'h991E: data = 8'b00000000;
            16'h991F: data = 8'b00000000;
            // code x992 (2-TH)
            16'h9920: data = 8'b00000000;
            16'h9921: data = 8'b00000000;
            16'h9922: data = 8'b10000000;
            16'h9923: data = 8'b10000000;
            16'h9924: data = 8'b10000000;
            16'h9925: data = 8'b10010100;
            16'h9926: data = 8'b10101010;
            16'h9927: data = 8'b10110010;
            16'h9928: data = 8'b10101010;
            16'h9929: data = 8'b10010010;
            16'h992A: data = 8'b11000110;
            16'h992B: data = 8'b01111100;
            16'h992C: data = 8'b00000000;
            16'h992D: data = 8'b00000000;
            16'h992E: data = 8'b00000000;
            16'h992F: data = 8'b00000000;
            // code x993 (3-TH)
            16'h9930: data = 8'b00000000;
            16'h9931: data = 8'b00000000;
            16'h9932: data = 8'b00000000;
            16'h9933: data = 8'b00000000;
            16'h9934: data = 8'b00000000;
            16'h9935: data = 8'b01101100;
            16'h9936: data = 8'b10010010;
            16'h9937: data = 8'b10010010;
            16'h9938: data = 8'b10000010;
            16'h9939: data = 8'b10100010;
            16'h993A: data = 8'b11010010;
            16'h993B: data = 8'b01100100;
            16'h993C: data = 8'b00000000;
            16'h993D: data = 8'b00000000;
            16'h993E: data = 8'b00000000;
            16'h993F: data = 8'b00000000;
            // code x994 (4-TH)
            16'h9940: data = 8'b00000000;
            16'h9941: data = 8'b00000000;
            16'h9942: data = 8'b00000010;
            16'h9943: data = 8'b00000010;
            16'h9944: data = 8'b00000100;
            16'h9945: data = 8'b01111000;
            16'h9946: data = 8'b11000000;
            16'h9947: data = 8'b10001000;
            16'h9948: data = 8'b10010100;
            16'h9949: data = 8'b10001100;
            16'h994A: data = 8'b11000010;
            16'h994B: data = 8'b01111110;
            16'h994C: data = 8'b00000000;
            16'h994D: data = 8'b00000000;
            16'h994E: data = 8'b00000000;
            16'h994F: data = 8'b00000000;
            // code x995 (5-TH)
            16'h9950: data = 8'b00000000;
            16'h9951: data = 8'b00000000;
            16'h9952: data = 8'b00000010;
            16'h9953: data = 8'b00100010;
            16'h9954: data = 8'b01010100;
            16'h9955: data = 8'b01111000;
            16'h9956: data = 8'b11000000;
            16'h9957: data = 8'b10001000;
            16'h9958: data = 8'b10010100;
            16'h9959: data = 8'b10001100;
            16'h995A: data = 8'b11000010;
            16'h995B: data = 8'b01111110;
            16'h995C: data = 8'b00000000;
            16'h995D: data = 8'b00000000;
            16'h995E: data = 8'b00000000;
            16'h995F: data = 8'b00000000;
            // code x996 (6-TH)
            16'h9960: data = 8'b00000000;
            16'h9961: data = 8'b00000000;
            16'h9962: data = 8'b10000000;
            16'h9963: data = 8'b11000000;
            16'h9964: data = 8'b01100000;
            16'h9965: data = 8'b00111000;
            16'h9966: data = 8'b00001100;
            16'h9967: data = 8'b01000110;
            16'h9968: data = 8'b10100010;
            16'h9969: data = 8'b11000010;
            16'h996A: data = 8'b10000110;
            16'h996B: data = 8'b01111100;
            16'h996C: data = 8'b00000000;
            16'h996D: data = 8'b00000000;
            16'h996E: data = 8'b00000000;
            16'h996F: data = 8'b00000000;
            // code x997 (7-TH)
            16'h9970: data = 8'b00000000;
            16'h9971: data = 8'b00000000;
            16'h9972: data = 8'b00000010;
            16'h9973: data = 8'b00000010;
            16'h9974: data = 8'b00000010;
            16'h9975: data = 8'b01101110;
            16'h9976: data = 8'b11010110;
            16'h9977: data = 8'b10010010;
            16'h9978: data = 8'b10010010;
            16'h9979: data = 8'b10100010;
            16'h997A: data = 8'b11010110;
            16'h997B: data = 8'b01101100;
            16'h997C: data = 8'b00000000;
            16'h997D: data = 8'b00000000;
            16'h997E: data = 8'b00000000;
            16'h997F: data = 8'b00000000;
            // code x998 (8-TH)
            16'h9980: data = 8'b00000000;
            16'h9981: data = 8'b00000000;
            16'h9982: data = 8'b00000010;
            16'h9983: data = 8'b00000010;
            16'h9984: data = 8'b00000010;
            16'h9985: data = 8'b00111110;
            16'h9986: data = 8'b01100000;
            16'h9987: data = 8'b11001100;
            16'h9988: data = 8'b10001010;
            16'h9989: data = 8'b10100110;
            16'h998A: data = 8'b10100110;
            16'h998B: data = 8'b01011100;
            16'h998C: data = 8'b00000000;
            16'h998D: data = 8'b00000000;
            16'h998E: data = 8'b00000000;
            16'h998F: data = 8'b00000000;
            // code x999 (9-TH)
            16'h9990: data = 8'b00000000;
            16'h9991: data = 8'b00000000;
            16'h9992: data = 8'b00000000;
            16'h9993: data = 8'b00000010;
            16'h9994: data = 8'b00000010;
            16'h9995: data = 8'b00111010;
            16'h9996: data = 8'b11101010;
            16'h9997: data = 8'b10100110;
            16'h9998: data = 8'b10010010;
            16'h9999: data = 8'b11101000;
            16'h999A: data = 8'b11010100;
            16'h999B: data = 8'b01100000;
            16'h999C: data = 8'b00000000;
            16'h999D: data = 8'b00000000;
            16'h999E: data = 8'b00000000;
            16'h999F: data = 8'b00000000;
			// default
			default: data = 8'b00000000;
		endcase
endmodule